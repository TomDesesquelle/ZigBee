
module FILTER ( Filter_In, CLK, RESET, ADC_Eocb, ADC_Convstb, ADC_Rdb, ADC_csb, 
        DAC_WRb, DAC_csb, LDACb, CLRb, Filter_Out );
  input [7:0] Filter_In;
  output [7:0] Filter_Out;
  input CLK, RESET, ADC_Eocb;
  output ADC_Convstb, ADC_Rdb, ADC_csb, DAC_WRb, DAC_csb, LDACb, CLRb;
  wire   ADC_Rdb, DAC_WRb, Delay_Line_sample_shift, Buff_OE, req_ADC2F,
         ack_F2ADC, req_F2DAC, \U1/n53 , \U1/n52 , \U1/n51 , \U1/n50 ,
         \U1/n49 , \U1/n48 , \U1/n47 , \U1/n46 , \U1/n45 , \U1/n44 , \U1/n43 ,
         \U1/n42 , \U1/n41 , \U1/n40 , \U1/n39 , \U1/n38 , \U1/n37 , \U1/n36 ,
         \U1/n35 , \U1/n34 , \U1/n33 , \U1/n32 , \U1/n31 , \U1/n30 , \U1/n29 ,
         \U1/n28 , \U1/n27 , \U1/n26 , \U1/n25 , \U1/n24 , \U1/n23 , \U1/n22 ,
         \U1/n21 , \U1/n20 , \U1/n19 , \U1/n18 , \U1/n17 , \U1/n16 , \U1/n15 ,
         \U1/n14 , \U1/n13 , \U1/n12 , \U1/n11 , \U1/n9 , \U1/n7 , \U1/n6 ,
         \U1/n5 , \U1/n4 , \U1/n3 , \U1/n2 , \U2/n741 , \U2/n740 , \U2/n739 ,
         \U2/n738 , \U2/n737 , \U2/n736 , \U2/n735 , \U2/n734 , \U2/n733 ,
         \U2/n732 , \U2/n731 , \U2/n730 , \U2/n729 , \U2/n728 , \U2/n727 ,
         \U2/n726 , \U2/n725 , \U2/n724 , \U2/n723 , \U2/n722 , \U2/n721 ,
         \U2/n720 , \U2/n719 , \U2/n718 , \U2/n717 , \U2/n716 , \U2/n715 ,
         \U2/n714 , \U2/n713 , \U2/n712 , \U2/n711 , \U2/n710 , \U2/n709 ,
         \U2/n708 , \U2/n707 , \U2/n706 , \U2/n705 , \U2/n704 , \U2/n703 ,
         \U2/n702 , \U2/n701 , \U2/n700 , \U2/n699 , \U2/n698 , \U2/n697 ,
         \U2/n696 , \U2/n695 , \U2/n694 , \U2/n693 , \U2/n692 , \U2/n691 ,
         \U2/n690 , \U2/n689 , \U2/n688 , \U2/n687 , \U2/n686 , \U2/n685 ,
         \U2/n684 , \U2/n683 , \U2/n682 , \U2/n681 , \U2/n680 , \U2/n679 ,
         \U2/n678 , \U2/n677 , \U2/n676 , \U2/n675 , \U2/n674 , \U2/n673 ,
         \U2/n672 , \U2/n671 , \U2/n670 , \U2/n669 , \U2/n668 , \U2/n667 ,
         \U2/n666 , \U2/n665 , \U2/n664 , \U2/n663 , \U2/n662 , \U2/n661 ,
         \U2/n660 , \U2/n659 , \U2/n658 , \U2/n657 , \U2/n656 , \U2/n655 ,
         \U2/n654 , \U2/n653 , \U2/n652 , \U2/n651 , \U2/n650 , \U2/n649 ,
         \U2/n648 , \U2/n647 , \U2/n646 , \U2/n645 , \U2/n644 , \U2/n643 ,
         \U2/n642 , \U2/n641 , \U2/n640 , \U2/n639 , \U2/n638 , \U2/n637 ,
         \U2/n636 , \U2/n635 , \U2/n634 , \U2/n633 , \U2/n632 , \U2/n631 ,
         \U2/n630 , \U2/n629 , \U2/n628 , \U2/n627 , \U2/n626 , \U2/n625 ,
         \U2/n624 , \U2/n623 , \U2/n622 , \U2/n621 , \U2/n620 , \U2/n619 ,
         \U2/n618 , \U2/n617 , \U2/n616 , \U2/n615 , \U2/n614 , \U2/n613 ,
         \U2/n612 , \U2/n611 , \U2/n610 , \U2/n609 , \U2/n608 , \U2/n607 ,
         \U2/n606 , \U2/n605 , \U2/n604 , \U2/n603 , \U2/n602 , \U2/n601 ,
         \U2/n600 , \U2/n599 , \U2/n598 , \U2/n597 , \U2/n596 , \U2/n595 ,
         \U2/n594 , \U2/n593 , \U2/n592 , \U2/n523 , \U2/n522 , \U2/n521 ,
         \U2/n520 , \U2/n519 , \U2/n518 , \U2/n517 , \U2/n516 , \U2/n391 ,
         \U2/n390 , \U2/n389 , \U2/n388 , \U2/n387 , \U2/n386 , \U2/n385 ,
         \U2/n384 , \U2/n383 , \U2/n382 , \U2/n381 , \U2/n380 , \U2/n379 ,
         \U2/n378 , \U2/n377 , \U2/n376 , \U2/n375 , \U2/n374 , \U2/n373 ,
         \U2/n372 , \U2/n371 , \U2/n370 , \U2/n369 , \U2/n368 , \U2/n367 ,
         \U2/n366 , \U2/n365 , \U2/n364 , \U2/n363 , \U2/n362 , \U2/n361 ,
         \U2/n360 , \U2/n359 , \U2/n358 , \U2/n357 , \U2/n356 , \U2/n355 ,
         \U2/n354 , \U2/n353 , \U2/n352 , \U2/n351 , \U2/n350 , \U2/n349 ,
         \U2/n348 , \U2/n347 , \U2/n346 , \U2/n345 , \U2/n344 , \U2/n343 ,
         \U2/n342 , \U2/n341 , \U2/n340 , \U2/n339 , \U2/n338 , \U2/n337 ,
         \U2/n336 , \U2/n335 , \U2/n334 , \U2/n333 , \U2/n332 , \U2/n331 ,
         \U2/n330 , \U2/n329 , \U2/n328 , \U2/n327 , \U2/n326 , \U2/n325 ,
         \U2/n324 , \U2/n323 , \U2/n322 , \U2/n321 , \U2/n320 , \U2/n319 ,
         \U2/n318 , \U2/n317 , \U2/n316 , \U2/n315 , \U2/n314 , \U2/n313 ,
         \U2/n312 , \U2/n311 , \U2/n310 , \U2/n309 , \U2/n308 , \U2/n307 ,
         \U2/n306 , \U2/n305 , \U2/n304 , \U2/n303 , \U2/n302 , \U2/n301 ,
         \U2/n300 , \U2/n299 , \U2/n298 , \U2/n297 , \U2/n296 , \U2/n295 ,
         \U2/n294 , \U2/n293 , \U2/n292 , \U2/n291 , \U2/n290 , \U2/n289 ,
         \U2/n288 , \U2/n287 , \U2/n286 , \U2/n285 , \U2/n284 , \U2/n280 ,
         \U2/n278 , \U2/n277 , \U2/n276 , \U2/n275 , \U2/n274 , \U2/n273 ,
         \U2/n272 , \U2/n271 , \U2/n270 , \U2/n269 , \U2/n268 , \U2/n267 ,
         \U2/n266 , \U2/n264 , \U2/n263 , \U2/n262 , \U2/n261 , \U2/n260 ,
         \U2/n259 , \U2/n258 , \U2/n257 , \U2/n256 , \U2/n255 , \U2/n254 ,
         \U2/n253 , \U2/n252 , \U2/n251 , \U2/n250 , \U2/n249 , \U2/n248 ,
         \U2/n247 , \U2/n246 , \U2/n245 , \U2/n244 , \U2/n243 , \U2/n242 ,
         \U2/n241 , \U2/n240 , \U2/n238 , \U2/n236 , \U2/n234 , \U2/n232 ,
         \U2/n230 , \U2/n228 , \U2/n226 , \U2/n32 , \U2/n31 , \U2/n30 ,
         \U2/n29 , \U2/n28 , \U2/n27 , \U2/n26 , \U2/n25 , \U2/n24 , \U2/n23 ,
         \U2/n22 , \U2/n21 , \U2/n20 , \U2/n19 , \U2/n18 , \U2/n17 , \U2/n16 ,
         \U2/n15 , \U2/n14 , \U2/n13 , \U2/n12 , \U2/n11 , \U2/n10 , \U2/n9 ,
         \U2/n8 , \U2/n7 , \U2/n6 , \U2/n5 , \U2/n4 , \U2/n3 , \U2/n2 ,
         \U2/n1 , \U2/n591 , \U2/n590 , \U2/n589 , \U2/n588 , \U2/n587 ,
         \U2/n586 , \U2/n585 , \U2/n584 , \U2/n583 , \U2/n582 , \U2/n581 ,
         \U2/n580 , \U2/n579 , \U2/n578 , \U2/n577 , \U2/n576 , \U2/n575 ,
         \U2/n574 , \U2/n573 , \U2/n572 , \U2/n571 , \U2/n570 , \U2/n569 ,
         \U2/n568 , \U2/n567 , \U2/n566 , \U2/n565 , \U2/n564 , \U2/n563 ,
         \U2/n562 , \U2/n561 , \U2/n560 , \U2/n559 , \U2/n558 , \U2/n557 ,
         \U2/n556 , \U2/n555 , \U2/n554 , \U2/n553 , \U2/n552 , \U2/n551 ,
         \U2/n550 , \U2/n549 , \U2/n548 , \U2/n547 , \U2/n546 , \U2/n545 ,
         \U2/n544 , \U2/n543 , \U2/n542 , \U2/n541 , \U2/n540 , \U2/n539 ,
         \U2/n538 , \U2/n537 , \U2/n536 , \U2/n535 , \U2/n534 , \U2/n533 ,
         \U2/n532 , \U2/n531 , \U2/n530 , \U2/n529 , \U2/n528 , \U2/n527 ,
         \U2/n526 , \U2/n525 , \U2/n524 , \U2/n515 , \U2/n514 , \U2/n513 ,
         \U2/n512 , \U2/n511 , \U2/n510 , \U2/n509 , \U2/n508 , \U2/n507 ,
         \U2/n506 , \U2/n505 , \U2/n504 , \U2/n503 , \U2/n502 , \U2/n501 ,
         \U2/n500 , \U2/n499 , \U2/n498 , \U2/n497 , \U2/n496 , \U2/n495 ,
         \U2/n494 , \U2/n493 , \U2/n492 , \U2/n491 , \U2/n490 , \U2/n489 ,
         \U2/n488 , \U2/n487 , \U2/n486 , \U2/n485 , \U2/n484 , \U2/n483 ,
         \U2/n482 , \U2/n481 , \U2/n480 , \U2/n479 , \U2/n478 , \U2/n477 ,
         \U2/n476 , \U2/n475 , \U2/n474 , \U2/n473 , \U2/n472 , \U2/n471 ,
         \U2/n470 , \U2/n469 , \U2/n468 , \U2/n467 , \U2/n466 , \U2/n465 ,
         \U2/n464 , \U2/n463 , \U2/n462 , \U2/n461 , \U2/n460 , \U2/n459 ,
         \U2/n458 , \U2/n457 , \U2/n456 , \U2/n455 , \U2/n454 , \U2/n453 ,
         \U2/n452 , \U2/n451 , \U2/n450 , \U2/n449 , \U2/n448 , \U2/n447 ,
         \U2/n446 , \U2/n445 , \U2/n444 , \U2/n443 , \U2/n442 , \U2/n441 ,
         \U2/n440 , \U2/n439 , \U2/n438 , \U2/n437 , \U2/n436 , \U2/n435 ,
         \U2/n434 , \U2/n433 , \U2/n432 , \U2/n431 , \U2/n430 , \U2/n429 ,
         \U2/n428 , \U2/n427 , \U2/n426 , \U2/n425 , \U2/n424 , \U2/n423 ,
         \U2/n422 , \U2/n421 , \U2/n420 , \U2/n419 , \U2/n418 , \U2/n417 ,
         \U2/n416 , \U2/n415 , \U2/n414 , \U2/n413 , \U2/n412 , \U2/n411 ,
         \U2/n410 , \U2/n409 , \U2/n408 , \U2/n407 , \U2/n406 , \U2/n405 ,
         \U2/n404 , \U2/n403 , \U2/n402 , \U2/n401 , \U2/n400 , \U2/n399 ,
         \U2/n398 , \U2/n397 , \U2/n396 , \U2/n395 , \U2/n394 , \U2/n393 ,
         \U2/n392 , \U2/x[0][7] , \U2/x[0][6] , \U2/x[0][5] , \U2/x[0][4] ,
         \U2/x[0][3] , \U2/x[0][2] , \U2/x[0][1] , \U2/x[0][0] , \U2/x[1][7] ,
         \U2/x[1][6] , \U2/x[1][5] , \U2/x[1][4] , \U2/x[1][3] , \U2/x[1][2] ,
         \U2/x[1][1] , \U2/x[1][0] , \U2/x[2][7] , \U2/x[2][6] , \U2/x[2][5] ,
         \U2/x[2][4] , \U2/x[2][3] , \U2/x[2][2] , \U2/x[2][1] , \U2/x[2][0] ,
         \U2/x[3][7] , \U2/x[3][6] , \U2/x[3][5] , \U2/x[3][4] , \U2/x[3][3] ,
         \U2/x[3][2] , \U2/x[3][1] , \U2/x[3][0] , \U2/x[8][7] , \U2/x[8][6] ,
         \U2/x[8][5] , \U2/x[8][4] , \U2/x[8][3] , \U2/x[8][2] , \U2/x[8][1] ,
         \U2/x[8][0] , \U2/x[9][7] , \U2/x[9][6] , \U2/x[9][5] , \U2/x[9][4] ,
         \U2/x[9][3] , \U2/x[9][2] , \U2/x[9][1] , \U2/x[9][0] , \U2/x[10][7] ,
         \U2/x[10][6] , \U2/x[10][5] , \U2/x[10][4] , \U2/x[10][3] ,
         \U2/x[10][2] , \U2/x[10][1] , \U2/x[10][0] , \U2/x[11][7] ,
         \U2/x[11][6] , \U2/x[11][5] , \U2/x[11][4] , \U2/x[11][3] ,
         \U2/x[11][2] , \U2/x[11][1] , \U2/x[11][0] , \U2/x[12][7] ,
         \U2/x[12][6] , \U2/x[12][5] , \U2/x[12][4] , \U2/x[12][3] ,
         \U2/x[12][2] , \U2/x[12][1] , \U2/x[12][0] , \U2/x[13][7] ,
         \U2/x[13][6] , \U2/x[13][5] , \U2/x[13][4] , \U2/x[13][3] ,
         \U2/x[13][2] , \U2/x[13][1] , \U2/x[13][0] , \U2/x[14][7] ,
         \U2/x[14][6] , \U2/x[14][5] , \U2/x[14][4] , \U2/x[14][3] ,
         \U2/x[14][2] , \U2/x[14][1] , \U2/x[14][0] , \U2/x[15][7] ,
         \U2/x[15][6] , \U2/x[15][5] , \U2/x[15][4] , \U2/x[15][3] ,
         \U2/x[15][2] , \U2/x[15][1] , \U2/x[15][0] , \U2/x[16][7] ,
         \U2/x[16][6] , \U2/x[16][5] , \U2/x[16][4] , \U2/x[16][3] ,
         \U2/x[16][2] , \U2/x[16][1] , \U2/x[16][0] , \U2/x[17][7] ,
         \U2/x[17][6] , \U2/x[17][5] , \U2/x[17][4] , \U2/x[17][3] ,
         \U2/x[17][2] , \U2/x[17][1] , \U2/x[17][0] , \U2/x[18][7] ,
         \U2/x[18][6] , \U2/x[18][5] , \U2/x[18][4] , \U2/x[18][3] ,
         \U2/x[18][2] , \U2/x[18][1] , \U2/x[18][0] , \U2/x[19][7] ,
         \U2/x[19][6] , \U2/x[19][5] , \U2/x[19][4] , \U2/x[19][3] ,
         \U2/x[19][2] , \U2/x[19][1] , \U2/x[19][0] , \U2/x[24][7] ,
         \U2/x[24][6] , \U2/x[24][5] , \U2/x[24][4] , \U2/x[24][3] ,
         \U2/x[24][2] , \U2/x[24][1] , \U2/x[24][0] , \U2/x[25][7] ,
         \U2/x[25][6] , \U2/x[25][5] , \U2/x[25][4] , \U2/x[25][3] ,
         \U2/x[25][2] , \U2/x[25][1] , \U2/x[25][0] , \U2/x[26][7] ,
         \U2/x[26][6] , \U2/x[26][5] , \U2/x[26][4] , \U2/x[26][3] ,
         \U2/x[26][2] , \U2/x[26][1] , \U2/x[26][0] , \U2/x[27][7] ,
         \U2/x[27][6] , \U2/x[27][5] , \U2/x[27][4] , \U2/x[27][3] ,
         \U2/x[27][2] , \U2/x[27][1] , \U2/x[27][0] , \U2/x[28][7] ,
         \U2/x[28][6] , \U2/x[28][5] , \U2/x[28][4] , \U2/x[28][3] ,
         \U2/x[28][2] , \U2/x[28][1] , \U2/x[28][0] , \U2/x[29][7] ,
         \U2/x[29][6] , \U2/x[29][5] , \U2/x[29][4] , \U2/x[29][3] ,
         \U2/x[29][2] , \U2/x[29][1] , \U2/x[29][0] , \U2/x[30][7] ,
         \U2/x[30][6] , \U2/x[30][5] , \U2/x[30][4] , \U2/x[30][3] ,
         \U2/x[30][2] , \U2/x[30][1] , \U2/x[30][0] , \U2/x[31][7] ,
         \U2/x[31][6] , \U2/x[31][5] , \U2/x[31][4] , \U2/x[31][3] ,
         \U2/x[31][2] , \U2/x[31][1] , \U2/x[31][0] , \U4/n42 , \U4/n41 ,
         \U4/n40 , \U4/n39 , \U4/n38 , \U4/n37 , \U4/n36 , \U4/n35 , \U4/n34 ,
         \U4/n33 , \U4/n32 , \U4/n31 , \U4/n30 , \U4/n29 , \U4/n28 , \U4/N49 ,
         \U4/N50 , \U4/N51 , \U4/N52 , \U4/N53 , \U4/N54 , \U4/N55 , \U4/N56 ,
         \U4/N57 , \U4/N58 , \U4/N59 , \U4/N60 , \U4/N61 , \U4/N62 , \U4/N63 ,
         \U4/N64 , \U4/N65 , \U4/N66 , \U4/N46 , \U4/N45 , \U4/N44 , \U4/N43 ,
         \U4/N42 , \U4/N41 , \U4/N40 , \U4/N39 , \U4/N38 , \U4/N37 , \U4/N36 ,
         \U4/N35 , \U4/N34 , \U4/N33 , \U4/N32 , \U4/N31 , \U4/N30 , \U4/N29 ,
         \U4/N28 , \U4/N27 , \U4/N21 , \U4/N20 , \U4/N19 , \U4/N18 , \U4/N17 ,
         \U4/N16 , \U4/N15 , \U4/N14 , \U4/N13 , \U4/N12 , \U4/N11 , \U4/N10 ,
         \U4/N9 , \U4/N8 , \U4/N7 , \U4/Accu_out[0] , \U4/Accu_out[1] ,
         \U4/Accu_out[2] , \U4/Accu_out[3] , \U4/Accu_out[4] ,
         \U4/Accu_out[5] , \U4/Accu_out[6] , \U4/Accu_out[7] ,
         \U4/Accu_out[8] , \U4/Accu_out[9] , \U4/Accu_out[10] ,
         \U4/Accu_out[11] , \U5/n11 , \U5/n10 , \U5/n9 , \U5/n8 , \U5/n7 ,
         \U5/n6 , \U5/n5 , \U5/n4 , \U5/n3 , \U5/n2 , \U5/n1 , \U5/n27 ,
         \U5/n26 , \U5/n25 , \U5/n24 , \U5/n23 , \U5/n22 , \U5/n21 , \U5/n20 ,
         \U5/n19 , \U5/n18 , \U5/n17 , \U5/n16 , \U5/n15 , \U5/n14 , \U5/n13 ,
         \U5/n12 , \U6/n50 , \U6/n48 , \U6/n47 , \U6/n46 , \U6/n44 , \U6/n43 ,
         \U6/n36 , \U6/n35 , \U6/n34 , \U6/n32 , \U6/n31 , \U6/n29 , \U6/n28 ,
         \U6/n27 , \U6/n26 , \U6/n25 , \U6/n24 , \U6/n23 , \U6/n16 , \U6/n13 ,
         \U6/n11 , \U6/n10 , \U6/n8 , \U6/n7 , \U6/n33 , \U6/n4 , \U6/n2 ,
         \U6/n42 , \U6/n41 , \U6/n40 , \U6/n39 , \U6/n38 , \U6/n37 , \U6/n14 ,
         \U7/n12 , \U7/n11 , \U7/n10 , \U7/n1 , \U7/n9 , \U7/n2 , \U7/n15 ,
         \U7/n14 , \U7/n13 , \U8/n5 , \U8/n1 , \U8/N5 , \U8/pre_req_F2DAC ,
         \U8/current_state , \U9/n11 , \U9/n10 , \U9/n9 , \U9/n8 , \U9/n7 ,
         \U9/n6 , \U9/n5 , \U9/n4 , \U9/n3 , \U9/n2 , \U9/n1 , \U9/n27 ,
         \U9/n26 , \U9/n25 , \U9/n24 , \U9/n23 , \U9/n22 , \U9/n21 , \U9/n20 ,
         \U9/n19 , \U9/n18 , \U9/n17 , \U9/n16 , \U9/n15 , \U9/n14 , \U9/n13 ,
         \U9/n12 , \U3/mult_19/n91 , \U3/mult_19/n90 , \U3/mult_19/n89 ,
         \U3/mult_19/n88 , \U3/mult_19/n87 , \U3/mult_19/n86 ,
         \U3/mult_19/n85 , \U3/mult_19/n84 , \U3/mult_19/n83 ,
         \U3/mult_19/n80 , \U3/mult_19/n79 , \U3/mult_19/n78 ,
         \U3/mult_19/n75 , \U3/mult_19/n72 , \U3/mult_19/n71 ,
         \U3/mult_19/n70 , \U3/mult_19/n67 , \U3/mult_19/n66 ,
         \U3/mult_19/n65 , \U3/mult_19/n64 , \U3/mult_19/n63 ,
         \U3/mult_19/n62 , \U3/mult_19/n54 , \U3/mult_19/n51 ,
         \U3/mult_19/A2[7] , \U3/mult_19/A2[8] , \U3/mult_19/A2[9] ,
         \U3/mult_19/A2[10] , \U3/mult_19/A2[11] , \U3/mult_19/A2[12] ,
         \U3/mult_19/A1[7] , \U3/mult_19/A1[8] , \U3/mult_19/A1[9] ,
         \U3/mult_19/A1[10] , \U3/mult_19/A1[11] , \U3/mult_19/A1[12] ,
         \U3/mult_19/SUMB[1][1] , \U3/mult_19/SUMB[1][2] ,
         \U3/mult_19/SUMB[1][3] , \U3/mult_19/SUMB[1][4] ,
         \U3/mult_19/SUMB[1][5] , \U3/mult_19/SUMB[1][6] ,
         \U3/mult_19/SUMB[2][1] , \U3/mult_19/SUMB[2][2] ,
         \U3/mult_19/SUMB[2][3] , \U3/mult_19/SUMB[2][4] ,
         \U3/mult_19/SUMB[2][5] , \U3/mult_19/SUMB[2][6] ,
         \U3/mult_19/SUMB[3][1] , \U3/mult_19/SUMB[3][2] ,
         \U3/mult_19/SUMB[3][3] , \U3/mult_19/SUMB[3][4] ,
         \U3/mult_19/SUMB[3][5] , \U3/mult_19/SUMB[3][6] ,
         \U3/mult_19/SUMB[4][1] , \U3/mult_19/SUMB[4][2] ,
         \U3/mult_19/SUMB[4][3] , \U3/mult_19/SUMB[4][4] ,
         \U3/mult_19/SUMB[4][5] , \U3/mult_19/SUMB[4][6] ,
         \U3/mult_19/SUMB[5][1] , \U3/mult_19/SUMB[5][2] ,
         \U3/mult_19/SUMB[5][3] , \U3/mult_19/SUMB[5][4] ,
         \U3/mult_19/SUMB[5][5] , \U3/mult_19/SUMB[5][6] ,
         \U3/mult_19/SUMB[6][1] , \U3/mult_19/SUMB[6][2] ,
         \U3/mult_19/SUMB[6][3] , \U3/mult_19/SUMB[6][4] ,
         \U3/mult_19/SUMB[6][5] , \U3/mult_19/SUMB[6][6] ,
         \U3/mult_19/SUMB[7][1] , \U3/mult_19/SUMB[7][2] ,
         \U3/mult_19/SUMB[7][3] , \U3/mult_19/SUMB[7][4] ,
         \U3/mult_19/SUMB[7][5] , \U3/mult_19/SUMB[7][6] ,
         \U3/mult_19/CARRYB[1][0] , \U3/mult_19/CARRYB[1][1] ,
         \U3/mult_19/CARRYB[1][2] , \U3/mult_19/CARRYB[1][3] ,
         \U3/mult_19/CARRYB[1][4] , \U3/mult_19/CARRYB[1][5] ,
         \U3/mult_19/CARRYB[1][6] , \U3/mult_19/CARRYB[2][0] ,
         \U3/mult_19/CARRYB[2][1] , \U3/mult_19/CARRYB[2][2] ,
         \U3/mult_19/CARRYB[2][3] , \U3/mult_19/CARRYB[2][4] ,
         \U3/mult_19/CARRYB[2][5] , \U3/mult_19/CARRYB[2][6] ,
         \U3/mult_19/CARRYB[3][0] , \U3/mult_19/CARRYB[3][1] ,
         \U3/mult_19/CARRYB[3][2] , \U3/mult_19/CARRYB[3][3] ,
         \U3/mult_19/CARRYB[3][4] , \U3/mult_19/CARRYB[3][5] ,
         \U3/mult_19/CARRYB[3][6] , \U3/mult_19/CARRYB[4][0] ,
         \U3/mult_19/CARRYB[4][1] , \U3/mult_19/CARRYB[4][2] ,
         \U3/mult_19/CARRYB[4][3] , \U3/mult_19/CARRYB[4][4] ,
         \U3/mult_19/CARRYB[4][5] , \U3/mult_19/CARRYB[4][6] ,
         \U3/mult_19/CARRYB[5][0] , \U3/mult_19/CARRYB[5][1] ,
         \U3/mult_19/CARRYB[5][2] , \U3/mult_19/CARRYB[5][3] ,
         \U3/mult_19/CARRYB[5][4] , \U3/mult_19/CARRYB[5][5] ,
         \U3/mult_19/CARRYB[5][6] , \U3/mult_19/CARRYB[6][0] ,
         \U3/mult_19/CARRYB[6][1] , \U3/mult_19/CARRYB[6][2] ,
         \U3/mult_19/CARRYB[6][3] , \U3/mult_19/CARRYB[6][4] ,
         \U3/mult_19/CARRYB[6][5] , \U3/mult_19/CARRYB[6][6] ,
         \U3/mult_19/CARRYB[7][0] , \U3/mult_19/CARRYB[7][1] ,
         \U3/mult_19/CARRYB[7][2] , \U3/mult_19/CARRYB[7][3] ,
         \U3/mult_19/CARRYB[7][4] , \U3/mult_19/CARRYB[7][5] ,
         \U3/mult_19/CARRYB[7][6] , \U3/mult_19/ab[0][1] ,
         \U3/mult_19/ab[0][2] , \U3/mult_19/ab[0][3] , \U3/mult_19/ab[0][4] ,
         \U3/mult_19/ab[0][5] , \U3/mult_19/ab[0][6] , \U3/mult_19/ab[0][7] ,
         \U3/mult_19/ab[1][0] , \U3/mult_19/ab[1][1] , \U3/mult_19/ab[1][2] ,
         \U3/mult_19/ab[1][3] , \U3/mult_19/ab[1][4] , \U3/mult_19/ab[1][5] ,
         \U3/mult_19/ab[1][6] , \U3/mult_19/ab[1][7] , \U3/mult_19/ab[2][0] ,
         \U3/mult_19/ab[2][1] , \U3/mult_19/ab[2][2] , \U3/mult_19/ab[2][3] ,
         \U3/mult_19/ab[2][4] , \U3/mult_19/ab[2][5] , \U3/mult_19/ab[2][6] ,
         \U3/mult_19/ab[2][7] , \U3/mult_19/ab[3][0] , \U3/mult_19/ab[3][1] ,
         \U3/mult_19/ab[3][2] , \U3/mult_19/ab[3][3] , \U3/mult_19/ab[3][4] ,
         \U3/mult_19/ab[3][5] , \U3/mult_19/ab[3][6] , \U3/mult_19/ab[3][7] ,
         \U3/mult_19/ab[4][0] , \U3/mult_19/ab[4][1] , \U3/mult_19/ab[4][2] ,
         \U3/mult_19/ab[4][3] , \U3/mult_19/ab[4][4] , \U3/mult_19/ab[4][5] ,
         \U3/mult_19/ab[4][6] , \U3/mult_19/ab[4][7] , \U3/mult_19/ab[5][0] ,
         \U3/mult_19/ab[5][1] , \U3/mult_19/ab[5][2] , \U3/mult_19/ab[5][3] ,
         \U3/mult_19/ab[5][4] , \U3/mult_19/ab[5][5] , \U3/mult_19/ab[5][6] ,
         \U3/mult_19/ab[5][7] , \U3/mult_19/ab[6][0] , \U3/mult_19/ab[6][1] ,
         \U3/mult_19/ab[6][2] , \U3/mult_19/ab[6][3] , \U3/mult_19/ab[6][4] ,
         \U3/mult_19/ab[6][5] , \U3/mult_19/ab[6][6] , \U3/mult_19/ab[6][7] ,
         \U3/mult_19/ab[7][0] , \U3/mult_19/ab[7][1] , \U3/mult_19/ab[7][2] ,
         \U3/mult_19/ab[7][3] , \U3/mult_19/ab[7][4] , \U3/mult_19/ab[7][5] ,
         \U3/mult_19/ab[7][6] , \U3/mult_19/ab[7][7] , \U4/add_27_aco/n20 ,
         \U4/add_27_aco/n18 , \U4/add_27_aco/n14 ,
         \U4/mult_add_27_aco/PROD_not[0] , \U4/mult_add_27_aco/PROD_not[1] ,
         \U4/mult_add_27_aco/PROD_not[2] , \U4/mult_add_27_aco/PROD_not[3] ,
         \U4/mult_add_27_aco/PROD_not[4] , \U4/mult_add_27_aco/PROD_not[5] ,
         \U4/mult_add_27_aco/PROD_not[6] , \U4/mult_add_27_aco/PROD_not[7] ,
         \U4/mult_add_27_aco/PROD_not[8] , \U4/mult_add_27_aco/PROD_not[9] ,
         \U4/mult_add_27_aco/PROD_not[10] , \U4/mult_add_27_aco/PROD_not[11] ,
         \U4/mult_add_27_aco/PROD_not[12] , \U4/mult_add_27_aco/PROD_not[14] ,
         \U4/mult_add_27_aco/PROD_not[15] , \U4/mult_add_27_aco/PROD_not[16] ,
         \U4/mult_add_27_aco/PROD_not[17] , \U4/mult_add_27_aco/PROD_not[18] ,
         \U4/mult_add_27_aco/PROD_not[19] , \U3/mult_19/FS_1/n39 ,
         \U3/mult_19/FS_1/n37 , \U3/mult_19/FS_1/n34 , \U3/mult_19/FS_1/n33 ,
         \U3/mult_19/FS_1/n32 , \U3/mult_19/FS_1/n31 , \U3/mult_19/FS_1/n29 ,
         \U3/mult_19/FS_1/n28 , \U3/mult_19/FS_1/n27 , \U3/mult_19/FS_1/n26 ,
         \U3/mult_19/FS_1/n25 , \U3/mult_19/FS_1/n24 , \U3/mult_19/FS_1/n23 ,
         \U3/mult_19/FS_1/n22 , \U3/mult_19/FS_1/n21 , \U3/mult_19/FS_1/n20 ,
         \U3/mult_19/FS_1/n19 , \U3/mult_19/FS_1/n18 , \U3/mult_19/FS_1/n17 ,
         \U3/mult_19/FS_1/n16 , \U3/mult_19/FS_1/n15 , \U3/mult_19/FS_1/n14 ,
         \U3/mult_19/FS_1/n13 , \U3/mult_19/FS_1/n12 , \U3/mult_19/FS_1/n11 ,
         \U3/mult_19/FS_1/n10 , \U3/mult_19/FS_1/n9 , n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263;
  wire   [4:0] Rom_Address;
  wire   [7:0] Rom_out;
  wire   [7:0] Filter_In_mem;
  wire   [7:0] Delay_Line_out;
  wire   [15:0] Mult_out;
  wire   [19:12] Accu_out;
  wire   [20:1] \U4/add_27_aco/carry ;
  assign ADC_csb = ADC_Rdb;
  assign DAC_csb = DAC_WRb;

  OAI212 \U1/U27  ( .A(Rom_Address[4]), .B(\U1/n48 ), .C(\U1/n49 ), .Q(
        Rom_out[1]) );
  OAI212 \U1/U26  ( .A(n232), .B(\U1/n29 ), .C(\U1/n7 ), .Q(\U1/n47 ) );
  OAI212 \U1/U25  ( .A(n233), .B(\U1/n12 ), .C(\U1/n47 ), .Q(\U1/n44 ) );
  OAI222 \U1/U14  ( .A(Rom_out[7]), .B(\U1/n36 ), .C(\U1/n37 ), .D(\U1/n38 ), 
        .Q(Rom_out[3]) );
  OAI212 \U1/U7  ( .A(\U1/n27 ), .B(\U1/n28 ), .C(\U1/n2 ), .Q(\U1/n21 ) );
  OAI222 \U2/U413  ( .A(n123), .B(\U2/n358 ), .C(n34), .D(\U2/n359 ), .Q(
        \U2/n692 ) );
  OAI222 \U2/U412  ( .A(n122), .B(\U2/n356 ), .C(n33), .D(n235), .Q(\U2/n693 )
         );
  OAI222 \U2/U399  ( .A(Rom_Address[4]), .B(\U2/n678 ), .C(\U2/n679 ), .D(
        \U1/n2 ), .Q(Delay_Line_out[1]) );
  OAI222 \U2/U376  ( .A(Rom_Address[4]), .B(\U2/n656 ), .C(\U2/n657 ), .D(
        \U1/n2 ), .Q(Delay_Line_out[2]) );
  OAI222 \U2/U353  ( .A(Rom_Address[4]), .B(\U2/n634 ), .C(\U2/n635 ), .D(
        \U1/n2 ), .Q(Delay_Line_out[3]) );
  OAI222 \U2/U344  ( .A(n139), .B(\U2/n358 ), .C(n51), .D(n236), .Q(\U2/n626 )
         );
  OAI222 \U2/U343  ( .A(n138), .B(\U2/n356 ), .C(n50), .D(n235), .Q(\U2/n627 )
         );
  OAI222 \U2/U333  ( .A(n137), .B(\U2/n358 ), .C(n49), .D(n236), .Q(\U2/n616 )
         );
  OAI222 \U2/U332  ( .A(n25), .B(\U2/n356 ), .C(n18), .D(n235), .Q(\U2/n617 )
         );
  OAI222 \U2/U321  ( .A(n136), .B(\U2/n358 ), .C(n48), .D(n236), .Q(\U2/n604 )
         );
  OAI222 \U2/U320  ( .A(n135), .B(\U2/n356 ), .C(n47), .D(\U2/n357 ), .Q(
        \U2/n605 ) );
  OAI222 \U2/U310  ( .A(n134), .B(\U2/n358 ), .C(n46), .D(n236), .Q(\U2/n594 )
         );
  OAI222 \U2/U309  ( .A(n24), .B(\U2/n356 ), .C(n17), .D(\U2/n357 ), .Q(
        \U2/n595 ) );
  OAI222 \U2/U298  ( .A(n147), .B(\U2/n358 ), .C(n29), .D(n236), .Q(\U2/n390 )
         );
  OAI222 \U2/U297  ( .A(n146), .B(\U2/n356 ), .C(n55), .D(\U2/n357 ), .Q(
        \U2/n391 ) );
  OAI222 \U2/U287  ( .A(n145), .B(\U2/n358 ), .C(n54), .D(n236), .Q(\U2/n380 )
         );
  OAI222 \U2/U286  ( .A(n144), .B(\U2/n356 ), .C(n28), .D(\U2/n357 ), .Q(
        \U2/n381 ) );
  OAI222 \U2/U284  ( .A(Rom_Address[4]), .B(\U2/n376 ), .C(\U2/n377 ), .D(
        \U1/n2 ), .Q(Delay_Line_out[6]) );
  OAI222 \U2/U275  ( .A(n143), .B(\U2/n358 ), .C(n27), .D(n236), .Q(\U2/n368 )
         );
  OAI222 \U2/U274  ( .A(n142), .B(\U2/n356 ), .C(n53), .D(\U2/n357 ), .Q(
        \U2/n369 ) );
  OAI222 \U2/U264  ( .A(n141), .B(\U2/n358 ), .C(n52), .D(n236), .Q(\U2/n354 )
         );
  OAI222 \U2/U263  ( .A(n140), .B(\U2/n356 ), .C(n26), .D(\U2/n357 ), .Q(
        \U2/n355 ) );
  OAI222 \U2/U226  ( .A(n238), .B(n216), .C(n251), .D(n67), .Q(\U2/n392 ) );
  OAI222 \U2/U225  ( .A(n239), .B(n215), .C(n251), .D(n66), .Q(\U2/n393 ) );
  OAI222 \U2/U224  ( .A(n240), .B(n222), .C(n251), .D(n120), .Q(\U2/n394 ) );
  OAI222 \U2/U223  ( .A(n239), .B(n221), .C(n251), .D(n119), .Q(\U2/n395 ) );
  OAI222 \U2/U222  ( .A(n240), .B(n220), .C(n251), .D(n118), .Q(\U2/n396 ) );
  OAI222 \U2/U221  ( .A(n241), .B(n219), .C(n251), .D(n117), .Q(\U2/n397 ) );
  OAI222 \U2/U220  ( .A(n244), .B(n218), .C(n252), .D(n116), .Q(\U2/n398 ) );
  OAI222 \U2/U219  ( .A(n244), .B(n217), .C(n252), .D(n115), .Q(\U2/n399 ) );
  OAI222 \U2/U218  ( .A(n241), .B(n67), .C(n252), .D(n159), .Q(\U2/n400 ) );
  OAI222 \U2/U217  ( .A(n242), .B(n66), .C(n252), .D(n158), .Q(\U2/n401 ) );
  OAI222 \U2/U216  ( .A(n241), .B(n120), .C(n252), .D(n206), .Q(\U2/n402 ) );
  OAI222 \U2/U215  ( .A(n242), .B(n119), .C(n252), .D(n205), .Q(\U2/n403 ) );
  OAI222 \U2/U214  ( .A(n244), .B(n118), .C(n253), .D(n204), .Q(\U2/n404 ) );
  OAI222 \U2/U213  ( .A(n244), .B(n117), .C(n253), .D(n203), .Q(\U2/n405 ) );
  OAI222 \U2/U212  ( .A(n243), .B(n116), .C(n253), .D(n202), .Q(\U2/n406 ) );
  OAI222 \U2/U211  ( .A(n240), .B(n115), .C(n253), .D(n201), .Q(\U2/n407 ) );
  OAI222 \U2/U210  ( .A(n237), .B(n159), .C(n253), .D(n65), .Q(\U2/n408 ) );
  OAI222 \U2/U209  ( .A(n238), .B(n158), .C(n253), .D(n64), .Q(\U2/n409 ) );
  OAI222 \U2/U208  ( .A(n240), .B(n206), .C(n254), .D(n114), .Q(\U2/n410 ) );
  OAI222 \U2/U207  ( .A(n238), .B(n205), .C(n254), .D(n113), .Q(\U2/n411 ) );
  OAI222 \U2/U206  ( .A(n240), .B(n204), .C(n254), .D(n112), .Q(\U2/n412 ) );
  OAI222 \U2/U205  ( .A(n241), .B(n203), .C(n254), .D(n111), .Q(\U2/n413 ) );
  OAI222 \U2/U204  ( .A(n242), .B(n202), .C(n254), .D(n110), .Q(\U2/n414 ) );
  OAI222 \U2/U203  ( .A(n242), .B(n201), .C(n254), .D(n109), .Q(\U2/n415 ) );
  OAI222 \U2/U202  ( .A(n243), .B(n65), .C(n251), .D(n21), .Q(\U2/n416 ) );
  OAI222 \U2/U201  ( .A(n243), .B(n64), .C(n252), .D(n20), .Q(\U2/n417 ) );
  OAI222 \U2/U200  ( .A(n244), .B(n114), .C(n253), .D(n22), .Q(\U2/n418 ) );
  OAI222 \U2/U199  ( .A(n244), .B(n113), .C(n254), .D(n23), .Q(\U2/n419 ) );
  OAI222 \U2/U198  ( .A(n244), .B(n112), .C(n253), .D(n25), .Q(\U2/n420 ) );
  OAI222 \U2/U197  ( .A(n243), .B(n111), .C(n254), .D(n24), .Q(\U2/n421 ) );
  OAI222 \U2/U196  ( .A(n242), .B(n110), .C(n255), .D(n144), .Q(\U2/n422 ) );
  OAI222 \U2/U195  ( .A(n242), .B(n109), .C(n255), .D(n140), .Q(\U2/n423 ) );
  OAI222 \U2/U194  ( .A(n241), .B(n21), .C(n255), .D(n16), .Q(\U2/n424 ) );
  OAI222 \U2/U193  ( .A(n243), .B(n20), .C(n255), .D(n124), .Q(\U2/n425 ) );
  OAI222 \U2/U192  ( .A(n239), .B(n22), .C(n255), .D(n41), .Q(\U2/n426 ) );
  OAI222 \U2/U191  ( .A(n240), .B(n23), .C(n255), .D(n45), .Q(\U2/n427 ) );
  OAI222 \U2/U190  ( .A(n243), .B(n25), .C(n253), .D(n18), .Q(\U2/n428 ) );
  OAI222 \U2/U189  ( .A(n244), .B(n24), .C(n252), .D(n17), .Q(\U2/n429 ) );
  OAI222 \U2/U188  ( .A(n240), .B(n144), .C(n255), .D(n28), .Q(\U2/n430 ) );
  OAI222 \U2/U187  ( .A(n237), .B(n140), .C(n256), .D(n26), .Q(\U2/n431 ) );
  OAI222 \U2/U186  ( .A(n242), .B(n16), .C(n255), .D(n127), .Q(\U2/n432 ) );
  OAI222 \U2/U185  ( .A(n238), .B(n124), .C(n256), .D(n15), .Q(\U2/n433 ) );
  OAI222 \U2/U184  ( .A(n241), .B(n41), .C(n256), .D(n130), .Q(\U2/n434 ) );
  OAI222 \U2/U183  ( .A(n240), .B(n45), .C(n256), .D(n133), .Q(\U2/n435 ) );
  OAI222 \U2/U182  ( .A(n242), .B(n18), .C(n256), .D(n137), .Q(\U2/n436 ) );
  OAI222 \U2/U181  ( .A(n239), .B(n17), .C(n256), .D(n134), .Q(\U2/n437 ) );
  OAI222 \U2/U180  ( .A(n241), .B(n28), .C(n256), .D(n145), .Q(\U2/n438 ) );
  OAI222 \U2/U179  ( .A(n237), .B(n26), .C(n256), .D(n141), .Q(\U2/n439 ) );
  OAI222 \U2/U178  ( .A(n242), .B(n127), .C(n251), .D(n37), .Q(\U2/n440 ) );
  OAI222 \U2/U177  ( .A(n241), .B(n15), .C(n252), .D(n32), .Q(\U2/n441 ) );
  OAI222 \U2/U176  ( .A(n244), .B(n130), .C(n257), .D(n40), .Q(\U2/n442 ) );
  OAI222 \U2/U175  ( .A(n241), .B(n133), .C(n258), .D(n44), .Q(\U2/n443 ) );
  OAI222 \U2/U174  ( .A(n242), .B(n137), .C(n257), .D(n49), .Q(\U2/n444 ) );
  OAI222 \U2/U173  ( .A(n243), .B(n134), .C(n258), .D(n46), .Q(\U2/n445 ) );
  OAI222 \U2/U172  ( .A(n244), .B(n145), .C(n257), .D(n54), .Q(\U2/n446 ) );
  OAI222 \U2/U171  ( .A(n243), .B(n141), .C(n257), .D(n52), .Q(\U2/n447 ) );
  OAI222 \U2/U170  ( .A(n243), .B(n37), .C(n257), .D(n157), .Q(\U2/n448 ) );
  OAI222 \U2/U169  ( .A(n239), .B(n32), .C(n257), .D(n156), .Q(\U2/n449 ) );
  OAI222 \U2/U168  ( .A(n240), .B(n40), .C(n257), .D(n200), .Q(\U2/n450 ) );
  OAI222 \U2/U167  ( .A(n241), .B(n44), .C(n257), .D(n199), .Q(\U2/n451 ) );
  OAI222 \U2/U166  ( .A(n244), .B(n49), .C(n258), .D(n198), .Q(\U2/n452 ) );
  OAI222 \U2/U165  ( .A(n239), .B(n46), .C(n258), .D(n197), .Q(\U2/n453 ) );
  OAI222 \U2/U164  ( .A(n238), .B(n54), .C(n258), .D(n196), .Q(\U2/n454 ) );
  OAI222 \U2/U163  ( .A(n242), .B(n52), .C(n258), .D(n195), .Q(\U2/n455 ) );
  OAI222 \U2/U162  ( .A(n243), .B(n157), .C(n258), .D(n63), .Q(\U2/n456 ) );
  OAI222 \U2/U161  ( .A(n243), .B(n156), .C(n258), .D(n62), .Q(\U2/n457 ) );
  OAI222 \U2/U160  ( .A(n241), .B(n200), .C(n255), .D(n108), .Q(\U2/n458 ) );
  OAI222 \U2/U159  ( .A(n238), .B(n199), .C(n251), .D(n107), .Q(\U2/n459 ) );
  OAI222 \U2/U158  ( .A(n239), .B(n198), .C(n259), .D(n106), .Q(\U2/n460 ) );
  OAI222 \U2/U157  ( .A(n240), .B(n197), .C(n254), .D(n105), .Q(\U2/n461 ) );
  OAI222 \U2/U156  ( .A(n238), .B(n196), .C(n259), .D(n104), .Q(\U2/n462 ) );
  OAI222 \U2/U155  ( .A(n239), .B(n195), .C(n259), .D(n103), .Q(\U2/n463 ) );
  OAI222 \U2/U154  ( .A(n238), .B(n63), .C(n259), .D(n155), .Q(\U2/n464 ) );
  OAI222 \U2/U153  ( .A(n244), .B(n62), .C(n259), .D(n154), .Q(\U2/n465 ) );
  OAI222 \U2/U152  ( .A(n244), .B(n108), .C(n259), .D(n194), .Q(\U2/n466 ) );
  OAI222 \U2/U151  ( .A(n238), .B(n107), .C(n259), .D(n193), .Q(\U2/n467 ) );
  OAI222 \U2/U150  ( .A(n241), .B(n106), .C(n259), .D(n192), .Q(\U2/n468 ) );
  OAI222 \U2/U149  ( .A(n239), .B(n105), .C(n259), .D(n191), .Q(\U2/n469 ) );
  OAI222 \U2/U148  ( .A(n243), .B(n104), .C(n259), .D(n190), .Q(\U2/n470 ) );
  OAI222 \U2/U147  ( .A(n244), .B(n103), .C(n251), .D(n189), .Q(\U2/n471 ) );
  OAI222 \U2/U146  ( .A(n237), .B(n155), .C(n259), .D(n61), .Q(\U2/n472 ) );
  OAI222 \U2/U145  ( .A(n237), .B(n154), .C(n258), .D(n60), .Q(\U2/n473 ) );
  OAI222 \U2/U144  ( .A(n237), .B(n194), .C(n252), .D(n102), .Q(\U2/n474 ) );
  OAI222 \U2/U143  ( .A(n237), .B(n193), .C(n253), .D(n101), .Q(\U2/n475 ) );
  OAI222 \U2/U142  ( .A(n237), .B(n192), .C(n260), .D(n100), .Q(\U2/n476 ) );
  OAI222 \U2/U141  ( .A(n238), .B(n191), .C(n251), .D(n99), .Q(\U2/n477 ) );
  OAI222 \U2/U140  ( .A(n238), .B(n190), .C(n252), .D(n98), .Q(\U2/n478 ) );
  OAI222 \U2/U139  ( .A(n238), .B(n189), .C(n259), .D(n97), .Q(\U2/n479 ) );
  OAI222 \U2/U138  ( .A(n238), .B(n61), .C(n254), .D(n188), .Q(\U2/n480 ) );
  OAI222 \U2/U137  ( .A(n238), .B(n60), .C(n251), .D(n187), .Q(\U2/n481 ) );
  OAI222 \U2/U136  ( .A(n237), .B(n102), .C(n254), .D(n186), .Q(\U2/n482 ) );
  OAI222 \U2/U135  ( .A(n237), .B(n101), .C(n257), .D(n185), .Q(\U2/n483 ) );
  OAI222 \U2/U134  ( .A(n238), .B(n100), .C(n258), .D(n184), .Q(\U2/n484 ) );
  OAI222 \U2/U133  ( .A(n239), .B(n99), .C(n259), .D(n183), .Q(\U2/n485 ) );
  OAI222 \U2/U132  ( .A(n240), .B(n98), .C(n260), .D(n182), .Q(\U2/n486 ) );
  OAI222 \U2/U131  ( .A(n238), .B(n97), .C(n257), .D(n181), .Q(\U2/n487 ) );
  OAI222 \U2/U130  ( .A(n237), .B(n188), .C(n255), .D(n96), .Q(\U2/n488 ) );
  OAI222 \U2/U129  ( .A(n238), .B(n187), .C(n256), .D(n95), .Q(\U2/n489 ) );
  OAI222 \U2/U128  ( .A(n239), .B(n186), .C(n257), .D(n94), .Q(\U2/n490 ) );
  OAI222 \U2/U127  ( .A(n240), .B(n185), .C(n258), .D(n93), .Q(\U2/n491 ) );
  OAI222 \U2/U126  ( .A(n239), .B(n184), .C(n253), .D(n92), .Q(\U2/n492 ) );
  OAI222 \U2/U125  ( .A(n239), .B(n183), .C(n254), .D(n91), .Q(\U2/n493 ) );
  OAI222 \U2/U124  ( .A(n239), .B(n182), .C(n258), .D(n90), .Q(\U2/n494 ) );
  OAI222 \U2/U123  ( .A(n239), .B(n181), .C(n253), .D(n89), .Q(\U2/n495 ) );
  OAI222 \U2/U122  ( .A(n239), .B(n96), .C(n254), .D(n180), .Q(\U2/n496 ) );
  OAI222 \U2/U121  ( .A(n240), .B(n95), .C(n251), .D(n153), .Q(\U2/n497 ) );
  OAI222 \U2/U120  ( .A(n240), .B(n94), .C(n252), .D(n179), .Q(\U2/n498 ) );
  OAI222 \U2/U119  ( .A(n240), .B(n93), .C(n255), .D(n178), .Q(\U2/n499 ) );
  OAI222 \U2/U118  ( .A(n240), .B(n92), .C(n252), .D(n177), .Q(\U2/n500 ) );
  OAI222 \U2/U117  ( .A(n240), .B(n91), .C(n255), .D(n176), .Q(\U2/n501 ) );
  OAI222 \U2/U116  ( .A(n238), .B(n90), .C(n256), .D(n175), .Q(\U2/n502 ) );
  OAI222 \U2/U115  ( .A(n241), .B(n89), .C(n257), .D(n174), .Q(\U2/n503 ) );
  OAI222 \U2/U114  ( .A(n238), .B(n180), .C(n258), .D(n88), .Q(\U2/n504 ) );
  OAI222 \U2/U113  ( .A(n242), .B(n153), .C(n253), .D(n59), .Q(\U2/n505 ) );
  OAI222 \U2/U112  ( .A(n242), .B(n179), .C(n260), .D(n87), .Q(\U2/n506 ) );
  OAI222 \U2/U111  ( .A(n237), .B(n178), .C(n260), .D(n86), .Q(\U2/n507 ) );
  OAI222 \U2/U110  ( .A(n239), .B(n177), .C(n260), .D(n85), .Q(\U2/n508 ) );
  OAI222 \U2/U109  ( .A(n244), .B(n176), .C(n260), .D(n84), .Q(\U2/n509 ) );
  OAI222 \U2/U108  ( .A(n244), .B(n175), .C(n260), .D(n83), .Q(\U2/n510 ) );
  OAI222 \U2/U107  ( .A(n237), .B(n174), .C(n260), .D(n82), .Q(\U2/n511 ) );
  OAI222 \U2/U106  ( .A(n243), .B(n88), .C(n257), .D(n173), .Q(\U2/n512 ) );
  OAI222 \U2/U105  ( .A(n243), .B(n59), .C(n259), .D(n152), .Q(\U2/n513 ) );
  OAI222 \U2/U104  ( .A(n238), .B(n87), .C(n258), .D(n172), .Q(\U2/n514 ) );
  OAI222 \U2/U103  ( .A(n237), .B(n86), .C(n259), .D(n171), .Q(\U2/n515 ) );
  OAI222 \U2/U94  ( .A(n238), .B(n85), .C(n251), .D(n170), .Q(\U2/n524 ) );
  OAI222 \U2/U93  ( .A(n244), .B(n84), .C(n253), .D(n169), .Q(\U2/n525 ) );
  OAI222 \U2/U92  ( .A(n239), .B(n83), .C(n254), .D(n168), .Q(\U2/n526 ) );
  OAI222 \U2/U91  ( .A(n243), .B(n82), .C(n257), .D(n167), .Q(\U2/n527 ) );
  OAI222 \U2/U90  ( .A(n240), .B(n173), .C(n258), .D(n81), .Q(\U2/n528 ) );
  OAI222 \U2/U89  ( .A(n240), .B(n152), .C(n252), .D(n58), .Q(\U2/n529 ) );
  OAI222 \U2/U88  ( .A(n242), .B(n172), .C(n253), .D(n80), .Q(\U2/n530 ) );
  OAI222 \U2/U87  ( .A(n240), .B(n171), .C(n258), .D(n79), .Q(\U2/n531 ) );
  OAI222 \U2/U86  ( .A(n243), .B(n170), .C(n253), .D(n78), .Q(\U2/n532 ) );
  OAI222 \U2/U85  ( .A(n242), .B(n169), .C(n253), .D(n77), .Q(\U2/n533 ) );
  OAI222 \U2/U84  ( .A(n238), .B(n168), .C(n253), .D(n76), .Q(\U2/n534 ) );
  OAI222 \U2/U83  ( .A(n240), .B(n167), .C(n254), .D(n75), .Q(\U2/n535 ) );
  OAI222 \U2/U82  ( .A(n242), .B(n81), .C(n259), .D(n166), .Q(\U2/n536 ) );
  OAI222 \U2/U81  ( .A(n237), .B(n58), .C(n254), .D(n151), .Q(\U2/n537 ) );
  OAI222 \U2/U80  ( .A(n238), .B(n80), .C(n260), .D(n165), .Q(\U2/n538 ) );
  OAI222 \U2/U79  ( .A(n241), .B(n79), .C(n260), .D(n164), .Q(\U2/n539 ) );
  OAI222 \U2/U78  ( .A(n241), .B(n78), .C(n253), .D(n163), .Q(\U2/n540 ) );
  OAI222 \U2/U77  ( .A(n241), .B(n77), .C(n260), .D(n162), .Q(\U2/n541 ) );
  OAI222 \U2/U76  ( .A(n241), .B(n76), .C(n252), .D(n161), .Q(\U2/n542 ) );
  OAI222 \U2/U75  ( .A(n241), .B(n75), .C(n258), .D(n160), .Q(\U2/n543 ) );
  OAI222 \U2/U74  ( .A(n241), .B(n166), .C(n255), .D(n74), .Q(\U2/n544 ) );
  OAI222 \U2/U73  ( .A(n242), .B(n151), .C(n254), .D(n57), .Q(\U2/n545 ) );
  OAI222 \U2/U72  ( .A(n242), .B(n165), .C(n260), .D(n73), .Q(\U2/n546 ) );
  OAI222 \U2/U71  ( .A(n242), .B(n164), .C(n255), .D(n72), .Q(\U2/n547 ) );
  OAI222 \U2/U70  ( .A(n242), .B(n163), .C(n256), .D(n71), .Q(\U2/n548 ) );
  OAI222 \U2/U69  ( .A(n242), .B(n162), .C(n260), .D(n70), .Q(\U2/n549 ) );
  OAI222 \U2/U68  ( .A(n243), .B(n161), .C(n256), .D(n69), .Q(\U2/n550 ) );
  OAI222 \U2/U67  ( .A(n243), .B(n160), .C(n257), .D(n68), .Q(\U2/n551 ) );
  OAI222 \U2/U66  ( .A(n243), .B(n74), .C(n258), .D(n126), .Q(\U2/n552 ) );
  OAI222 \U2/U65  ( .A(n243), .B(n57), .C(n259), .D(n122), .Q(\U2/n553 ) );
  OAI222 \U2/U64  ( .A(n243), .B(n73), .C(n256), .D(n129), .Q(\U2/n554 ) );
  OAI222 \U2/U63  ( .A(n239), .B(n72), .C(n255), .D(n132), .Q(\U2/n555 ) );
  OAI222 \U2/U62  ( .A(n239), .B(n71), .C(n255), .D(n138), .Q(\U2/n556 ) );
  OAI222 \U2/U61  ( .A(n237), .B(n70), .C(n256), .D(n135), .Q(\U2/n557 ) );
  OAI222 \U2/U60  ( .A(n238), .B(n69), .C(n260), .D(n146), .Q(\U2/n558 ) );
  OAI222 \U2/U59  ( .A(n237), .B(n68), .C(n256), .D(n142), .Q(\U2/n559 ) );
  OAI222 \U2/U58  ( .A(n244), .B(n126), .C(n256), .D(n36), .Q(\U2/n560 ) );
  OAI222 \U2/U57  ( .A(n244), .B(n122), .C(n259), .D(n33), .Q(\U2/n561 ) );
  OAI222 \U2/U56  ( .A(n244), .B(n129), .C(n251), .D(n39), .Q(\U2/n562 ) );
  OAI222 \U2/U55  ( .A(n244), .B(n132), .C(n251), .D(n43), .Q(\U2/n563 ) );
  OAI222 \U2/U54  ( .A(n244), .B(n138), .C(n256), .D(n50), .Q(\U2/n564 ) );
  OAI222 \U2/U53  ( .A(n237), .B(n135), .C(n254), .D(n47), .Q(\U2/n565 ) );
  OAI222 \U2/U52  ( .A(n243), .B(n146), .C(n260), .D(n55), .Q(\U2/n566 ) );
  OAI222 \U2/U51  ( .A(n237), .B(n142), .C(n252), .D(n53), .Q(\U2/n567 ) );
  OAI222 \U2/U50  ( .A(n241), .B(n36), .C(n252), .D(n125), .Q(\U2/n568 ) );
  OAI222 \U2/U49  ( .A(n242), .B(n33), .C(n251), .D(n123), .Q(\U2/n569 ) );
  OAI222 \U2/U48  ( .A(n239), .B(n39), .C(n251), .D(n128), .Q(\U2/n570 ) );
  OAI222 \U2/U47  ( .A(n240), .B(n43), .C(n257), .D(n131), .Q(\U2/n571 ) );
  OAI222 \U2/U46  ( .A(n237), .B(n50), .C(n254), .D(n139), .Q(\U2/n572 ) );
  OAI222 \U2/U45  ( .A(n237), .B(n47), .C(n257), .D(n136), .Q(\U2/n573 ) );
  OAI222 \U2/U44  ( .A(n239), .B(n55), .C(n255), .D(n147), .Q(\U2/n574 ) );
  OAI222 \U2/U43  ( .A(n242), .B(n53), .C(n256), .D(n143), .Q(\U2/n575 ) );
  OAI222 \U2/U42  ( .A(n244), .B(n125), .C(n257), .D(n35), .Q(\U2/n576 ) );
  OAI222 \U2/U41  ( .A(n241), .B(n123), .C(n258), .D(n34), .Q(\U2/n577 ) );
  OAI222 \U2/U40  ( .A(n242), .B(n128), .C(n259), .D(n38), .Q(\U2/n578 ) );
  OAI222 \U2/U39  ( .A(n244), .B(n131), .C(n251), .D(n42), .Q(\U2/n579 ) );
  OAI222 \U2/U38  ( .A(n239), .B(n139), .C(n260), .D(n51), .Q(\U2/n580 ) );
  OAI222 \U2/U37  ( .A(n240), .B(n136), .C(n254), .D(n48), .Q(\U2/n581 ) );
  OAI222 \U2/U36  ( .A(n241), .B(n147), .C(n259), .D(n29), .Q(\U2/n582 ) );
  OAI222 \U2/U35  ( .A(n237), .B(n143), .C(n260), .D(n27), .Q(\U2/n583 ) );
  OAI222 \U2/U34  ( .A(n243), .B(n35), .C(n253), .D(n208), .Q(\U2/n584 ) );
  OAI222 \U2/U33  ( .A(n239), .B(n34), .C(n252), .D(n207), .Q(\U2/n585 ) );
  OAI222 \U2/U32  ( .A(n237), .B(n38), .C(n252), .D(n214), .Q(\U2/n586 ) );
  OAI222 \U2/U31  ( .A(n240), .B(n42), .C(n260), .D(n213), .Q(\U2/n587 ) );
  OAI222 \U2/U30  ( .A(n241), .B(n51), .C(n255), .D(n212), .Q(\U2/n588 ) );
  OAI222 \U2/U29  ( .A(n241), .B(n48), .C(n260), .D(n211), .Q(\U2/n589 ) );
  OAI222 \U2/U28  ( .A(n243), .B(n29), .C(n257), .D(n210), .Q(\U2/n590 ) );
  OAI222 \U2/U27  ( .A(n237), .B(n27), .C(n260), .D(n209), .Q(\U2/n591 ) );
  DF3 \U2/x_reg[31][0]  ( .D(\U2/n264 ), .C(CLK), .Q(\U2/x[31][0] ) );
  DF3 \U2/x_reg[31][1]  ( .D(\U2/n263 ), .C(CLK), .Q(\U2/x[31][1] ) );
  DF3 \U2/x_reg[31][2]  ( .D(\U2/n262 ), .C(CLK), .Q(\U2/x[31][2] ) );
  DF3 \U2/x_reg[31][3]  ( .D(\U2/n261 ), .C(CLK), .Q(\U2/x[31][3] ) );
  DF3 \U2/x_reg[31][4]  ( .D(\U2/n260 ), .C(CLK), .Q(\U2/x[31][4] ) );
  DF3 \U2/x_reg[31][5]  ( .D(\U2/n259 ), .C(CLK), .Q(\U2/x[31][5] ) );
  DF3 \U2/x_reg[31][6]  ( .D(\U2/n258 ), .C(CLK), .Q(\U2/x[31][6] ) );
  DF3 \U2/x_reg[31][7]  ( .D(\U2/n257 ), .C(CLK), .Q(\U2/x[31][7] ) );
  DF3 \U2/x_reg[30][0]  ( .D(\U2/n256 ), .C(CLK), .Q(\U2/x[30][0] ) );
  DF3 \U2/x_reg[30][1]  ( .D(\U2/n255 ), .C(CLK), .Q(\U2/x[30][1] ) );
  DF3 \U2/x_reg[30][2]  ( .D(\U2/n254 ), .C(CLK), .Q(\U2/x[30][2] ) );
  DF3 \U2/x_reg[30][3]  ( .D(\U2/n253 ), .C(CLK), .Q(\U2/x[30][3] ) );
  DF3 \U2/x_reg[30][4]  ( .D(\U2/n252 ), .C(CLK), .Q(\U2/x[30][4] ) );
  DF3 \U2/x_reg[30][5]  ( .D(\U2/n251 ), .C(CLK), .Q(\U2/x[30][5] ) );
  DF3 \U2/x_reg[30][6]  ( .D(\U2/n250 ), .C(CLK), .Q(\U2/x[30][6] ) );
  DF3 \U2/x_reg[30][7]  ( .D(\U2/n249 ), .C(CLK), .Q(\U2/x[30][7] ) );
  DF3 \U2/x_reg[29][0]  ( .D(\U2/n248 ), .C(CLK), .Q(\U2/x[29][0] ) );
  DF3 \U2/x_reg[29][1]  ( .D(\U2/n247 ), .C(CLK), .Q(\U2/x[29][1] ) );
  DF3 \U2/x_reg[29][2]  ( .D(\U2/n246 ), .C(CLK), .Q(\U2/x[29][2] ) );
  DF3 \U2/x_reg[29][3]  ( .D(\U2/n245 ), .C(CLK), .Q(\U2/x[29][3] ) );
  DF3 \U2/x_reg[29][4]  ( .D(\U2/n244 ), .C(CLK), .Q(\U2/x[29][4] ) );
  DF3 \U2/x_reg[29][5]  ( .D(\U2/n243 ), .C(CLK), .Q(\U2/x[29][5] ) );
  DF3 \U2/x_reg[29][6]  ( .D(\U2/n242 ), .C(CLK), .Q(\U2/x[29][6] ) );
  DF3 \U2/x_reg[29][7]  ( .D(\U2/n241 ), .C(CLK), .Q(\U2/x[29][7] ) );
  DF3 \U2/x_reg[28][0]  ( .D(\U2/n240 ), .C(CLK), .Q(\U2/x[28][0] ) );
  DF3 \U2/x_reg[28][1]  ( .D(\U2/n238 ), .C(CLK), .Q(\U2/x[28][1] ) );
  DF3 \U2/x_reg[28][2]  ( .D(\U2/n236 ), .C(CLK), .Q(\U2/x[28][2] ) );
  DF3 \U2/x_reg[28][3]  ( .D(\U2/n234 ), .C(CLK), .Q(\U2/x[28][3] ) );
  DF3 \U2/x_reg[28][4]  ( .D(\U2/n232 ), .C(CLK), .Q(\U2/x[28][4] ) );
  DF3 \U2/x_reg[28][5]  ( .D(\U2/n230 ), .C(CLK), .Q(\U2/x[28][5] ) );
  DF3 \U2/x_reg[28][6]  ( .D(\U2/n228 ), .C(CLK), .Q(\U2/x[28][6] ) );
  DF3 \U2/x_reg[28][7]  ( .D(\U2/n226 ), .C(CLK), .Q(\U2/x[28][7] ) );
  DF3 \U2/x_reg[27][0]  ( .D(\U2/n392 ), .C(CLK), .Q(\U2/x[27][0] ), .QN(n216)
         );
  DF3 \U2/x_reg[27][1]  ( .D(\U2/n393 ), .C(CLK), .Q(\U2/x[27][1] ), .QN(n215)
         );
  DF3 \U2/x_reg[27][2]  ( .D(\U2/n394 ), .C(CLK), .Q(\U2/x[27][2] ), .QN(n222)
         );
  DF3 \U2/x_reg[27][3]  ( .D(\U2/n395 ), .C(CLK), .Q(\U2/x[27][3] ), .QN(n221)
         );
  DF3 \U2/x_reg[27][4]  ( .D(\U2/n396 ), .C(CLK), .Q(\U2/x[27][4] ), .QN(n220)
         );
  DF3 \U2/x_reg[27][5]  ( .D(\U2/n397 ), .C(CLK), .Q(\U2/x[27][5] ), .QN(n219)
         );
  DF3 \U2/x_reg[27][6]  ( .D(\U2/n398 ), .C(CLK), .Q(\U2/x[27][6] ), .QN(n218)
         );
  DF3 \U2/x_reg[27][7]  ( .D(\U2/n399 ), .C(CLK), .Q(\U2/x[27][7] ), .QN(n217)
         );
  DF3 \U2/x_reg[26][0]  ( .D(\U2/n400 ), .C(CLK), .Q(\U2/x[26][0] ), .QN(n67)
         );
  DF3 \U2/x_reg[26][1]  ( .D(\U2/n401 ), .C(CLK), .Q(\U2/x[26][1] ), .QN(n66)
         );
  DF3 \U2/x_reg[26][2]  ( .D(\U2/n402 ), .C(CLK), .Q(\U2/x[26][2] ), .QN(n120)
         );
  DF3 \U2/x_reg[26][3]  ( .D(\U2/n403 ), .C(CLK), .Q(\U2/x[26][3] ), .QN(n119)
         );
  DF3 \U2/x_reg[26][4]  ( .D(\U2/n404 ), .C(CLK), .Q(\U2/x[26][4] ), .QN(n118)
         );
  DF3 \U2/x_reg[26][5]  ( .D(\U2/n405 ), .C(CLK), .Q(\U2/x[26][5] ), .QN(n117)
         );
  DF3 \U2/x_reg[26][6]  ( .D(\U2/n406 ), .C(CLK), .Q(\U2/x[26][6] ), .QN(n116)
         );
  DF3 \U2/x_reg[26][7]  ( .D(\U2/n407 ), .C(CLK), .Q(\U2/x[26][7] ), .QN(n115)
         );
  DF3 \U2/x_reg[25][0]  ( .D(\U2/n408 ), .C(CLK), .Q(\U2/x[25][0] ), .QN(n159)
         );
  DF3 \U2/x_reg[25][1]  ( .D(\U2/n409 ), .C(CLK), .Q(\U2/x[25][1] ), .QN(n158)
         );
  DF3 \U2/x_reg[25][2]  ( .D(\U2/n410 ), .C(CLK), .Q(\U2/x[25][2] ), .QN(n206)
         );
  DF3 \U2/x_reg[25][3]  ( .D(\U2/n411 ), .C(CLK), .Q(\U2/x[25][3] ), .QN(n205)
         );
  DF3 \U2/x_reg[25][4]  ( .D(\U2/n412 ), .C(CLK), .Q(\U2/x[25][4] ), .QN(n204)
         );
  DF3 \U2/x_reg[25][5]  ( .D(\U2/n413 ), .C(CLK), .Q(\U2/x[25][5] ), .QN(n203)
         );
  DF3 \U2/x_reg[25][6]  ( .D(\U2/n414 ), .C(CLK), .Q(\U2/x[25][6] ), .QN(n202)
         );
  DF3 \U2/x_reg[25][7]  ( .D(\U2/n415 ), .C(CLK), .Q(\U2/x[25][7] ), .QN(n201)
         );
  DF3 \U2/x_reg[24][0]  ( .D(\U2/n416 ), .C(CLK), .Q(\U2/x[24][0] ), .QN(n65)
         );
  DF3 \U2/x_reg[24][1]  ( .D(\U2/n417 ), .C(CLK), .Q(\U2/x[24][1] ), .QN(n64)
         );
  DF3 \U2/x_reg[24][2]  ( .D(\U2/n418 ), .C(CLK), .Q(\U2/x[24][2] ), .QN(n114)
         );
  DF3 \U2/x_reg[24][3]  ( .D(\U2/n419 ), .C(CLK), .Q(\U2/x[24][3] ), .QN(n113)
         );
  DF3 \U2/x_reg[24][4]  ( .D(\U2/n420 ), .C(CLK), .Q(\U2/x[24][4] ), .QN(n112)
         );
  DF3 \U2/x_reg[24][5]  ( .D(\U2/n421 ), .C(CLK), .Q(\U2/x[24][5] ), .QN(n111)
         );
  DF3 \U2/x_reg[24][6]  ( .D(\U2/n422 ), .C(CLK), .Q(\U2/x[24][6] ), .QN(n110)
         );
  DF3 \U2/x_reg[24][7]  ( .D(\U2/n423 ), .C(CLK), .Q(\U2/x[24][7] ), .QN(n109)
         );
  DF3 \U2/x_reg[23][0]  ( .D(\U2/n424 ), .C(CLK), .QN(n21) );
  DF3 \U2/x_reg[23][1]  ( .D(\U2/n425 ), .C(CLK), .QN(n20) );
  DF3 \U2/x_reg[23][2]  ( .D(\U2/n426 ), .C(CLK), .QN(n22) );
  DF3 \U2/x_reg[23][3]  ( .D(\U2/n427 ), .C(CLK), .QN(n23) );
  DF3 \U2/x_reg[23][4]  ( .D(\U2/n428 ), .C(CLK), .QN(n25) );
  DF3 \U2/x_reg[23][5]  ( .D(\U2/n429 ), .C(CLK), .QN(n24) );
  DF3 \U2/x_reg[23][6]  ( .D(\U2/n430 ), .C(CLK), .QN(n144) );
  DF3 \U2/x_reg[23][7]  ( .D(\U2/n431 ), .C(CLK), .QN(n140) );
  DF3 \U2/x_reg[22][0]  ( .D(\U2/n432 ), .C(CLK), .QN(n16) );
  DF3 \U2/x_reg[22][1]  ( .D(\U2/n433 ), .C(CLK), .QN(n124) );
  DF3 \U2/x_reg[22][2]  ( .D(\U2/n434 ), .C(CLK), .QN(n41) );
  DF3 \U2/x_reg[22][3]  ( .D(\U2/n435 ), .C(CLK), .QN(n45) );
  DF3 \U2/x_reg[22][4]  ( .D(\U2/n436 ), .C(CLK), .QN(n18) );
  DF3 \U2/x_reg[22][5]  ( .D(\U2/n437 ), .C(CLK), .QN(n17) );
  DF3 \U2/x_reg[22][6]  ( .D(\U2/n438 ), .C(CLK), .QN(n28) );
  DF3 \U2/x_reg[22][7]  ( .D(\U2/n439 ), .C(CLK), .QN(n26) );
  DF3 \U2/x_reg[21][0]  ( .D(\U2/n440 ), .C(CLK), .QN(n127) );
  DF3 \U2/x_reg[21][1]  ( .D(\U2/n441 ), .C(CLK), .QN(n15) );
  DF3 \U2/x_reg[21][2]  ( .D(\U2/n442 ), .C(CLK), .QN(n130) );
  DF3 \U2/x_reg[21][3]  ( .D(\U2/n443 ), .C(CLK), .QN(n133) );
  DF3 \U2/x_reg[21][4]  ( .D(\U2/n444 ), .C(CLK), .QN(n137) );
  DF3 \U2/x_reg[21][5]  ( .D(\U2/n445 ), .C(CLK), .QN(n134) );
  DF3 \U2/x_reg[21][6]  ( .D(\U2/n446 ), .C(CLK), .QN(n145) );
  DF3 \U2/x_reg[21][7]  ( .D(\U2/n447 ), .C(CLK), .QN(n141) );
  DF3 \U2/x_reg[20][0]  ( .D(\U2/n448 ), .C(CLK), .QN(n37) );
  DF3 \U2/x_reg[20][1]  ( .D(\U2/n449 ), .C(CLK), .QN(n32) );
  DF3 \U2/x_reg[20][2]  ( .D(\U2/n450 ), .C(CLK), .QN(n40) );
  DF3 \U2/x_reg[20][3]  ( .D(\U2/n451 ), .C(CLK), .QN(n44) );
  DF3 \U2/x_reg[20][4]  ( .D(\U2/n452 ), .C(CLK), .QN(n49) );
  DF3 \U2/x_reg[20][5]  ( .D(\U2/n453 ), .C(CLK), .QN(n46) );
  DF3 \U2/x_reg[20][6]  ( .D(\U2/n454 ), .C(CLK), .QN(n54) );
  DF3 \U2/x_reg[20][7]  ( .D(\U2/n455 ), .C(CLK), .QN(n52) );
  DF3 \U2/x_reg[19][0]  ( .D(\U2/n456 ), .C(CLK), .Q(\U2/x[19][0] ), .QN(n157)
         );
  DF3 \U2/x_reg[19][1]  ( .D(\U2/n457 ), .C(CLK), .Q(\U2/x[19][1] ), .QN(n156)
         );
  DF3 \U2/x_reg[19][2]  ( .D(\U2/n458 ), .C(CLK), .Q(\U2/x[19][2] ), .QN(n200)
         );
  DF3 \U2/x_reg[19][3]  ( .D(\U2/n459 ), .C(CLK), .Q(\U2/x[19][3] ), .QN(n199)
         );
  DF3 \U2/x_reg[19][4]  ( .D(\U2/n460 ), .C(CLK), .Q(\U2/x[19][4] ), .QN(n198)
         );
  DF3 \U2/x_reg[19][5]  ( .D(\U2/n461 ), .C(CLK), .Q(\U2/x[19][5] ), .QN(n197)
         );
  DF3 \U2/x_reg[19][6]  ( .D(\U2/n462 ), .C(CLK), .Q(\U2/x[19][6] ), .QN(n196)
         );
  DF3 \U2/x_reg[19][7]  ( .D(\U2/n463 ), .C(CLK), .Q(\U2/x[19][7] ), .QN(n195)
         );
  DF3 \U2/x_reg[18][0]  ( .D(\U2/n464 ), .C(CLK), .Q(\U2/x[18][0] ), .QN(n63)
         );
  DF3 \U2/x_reg[18][1]  ( .D(\U2/n465 ), .C(CLK), .Q(\U2/x[18][1] ), .QN(n62)
         );
  DF3 \U2/x_reg[18][2]  ( .D(\U2/n466 ), .C(CLK), .Q(\U2/x[18][2] ), .QN(n108)
         );
  DF3 \U2/x_reg[18][3]  ( .D(\U2/n467 ), .C(CLK), .Q(\U2/x[18][3] ), .QN(n107)
         );
  DF3 \U2/x_reg[18][4]  ( .D(\U2/n468 ), .C(CLK), .Q(\U2/x[18][4] ), .QN(n106)
         );
  DF3 \U2/x_reg[18][5]  ( .D(\U2/n469 ), .C(CLK), .Q(\U2/x[18][5] ), .QN(n105)
         );
  DF3 \U2/x_reg[18][6]  ( .D(\U2/n470 ), .C(CLK), .Q(\U2/x[18][6] ), .QN(n104)
         );
  DF3 \U2/x_reg[18][7]  ( .D(\U2/n471 ), .C(CLK), .Q(\U2/x[18][7] ), .QN(n103)
         );
  DF3 \U2/x_reg[17][0]  ( .D(\U2/n472 ), .C(CLK), .Q(\U2/x[17][0] ), .QN(n155)
         );
  DF3 \U2/x_reg[17][1]  ( .D(\U2/n473 ), .C(CLK), .Q(\U2/x[17][1] ), .QN(n154)
         );
  DF3 \U2/x_reg[17][2]  ( .D(\U2/n474 ), .C(CLK), .Q(\U2/x[17][2] ), .QN(n194)
         );
  DF3 \U2/x_reg[17][3]  ( .D(\U2/n475 ), .C(CLK), .Q(\U2/x[17][3] ), .QN(n193)
         );
  DF3 \U2/x_reg[17][4]  ( .D(\U2/n476 ), .C(CLK), .Q(\U2/x[17][4] ), .QN(n192)
         );
  DF3 \U2/x_reg[17][5]  ( .D(\U2/n477 ), .C(CLK), .Q(\U2/x[17][5] ), .QN(n191)
         );
  DF3 \U2/x_reg[17][6]  ( .D(\U2/n478 ), .C(CLK), .Q(\U2/x[17][6] ), .QN(n190)
         );
  DF3 \U2/x_reg[17][7]  ( .D(\U2/n479 ), .C(CLK), .Q(\U2/x[17][7] ), .QN(n189)
         );
  DF3 \U2/x_reg[16][0]  ( .D(\U2/n480 ), .C(CLK), .Q(\U2/x[16][0] ), .QN(n61)
         );
  DF3 \U2/x_reg[16][1]  ( .D(\U2/n481 ), .C(CLK), .Q(\U2/x[16][1] ), .QN(n60)
         );
  DF3 \U2/x_reg[16][2]  ( .D(\U2/n482 ), .C(CLK), .Q(\U2/x[16][2] ), .QN(n102)
         );
  DF3 \U2/x_reg[16][3]  ( .D(\U2/n483 ), .C(CLK), .Q(\U2/x[16][3] ), .QN(n101)
         );
  DF3 \U2/x_reg[16][4]  ( .D(\U2/n484 ), .C(CLK), .Q(\U2/x[16][4] ), .QN(n100)
         );
  DF3 \U2/x_reg[16][5]  ( .D(\U2/n485 ), .C(CLK), .Q(\U2/x[16][5] ), .QN(n99)
         );
  DF3 \U2/x_reg[16][6]  ( .D(\U2/n486 ), .C(CLK), .Q(\U2/x[16][6] ), .QN(n98)
         );
  DF3 \U2/x_reg[16][7]  ( .D(\U2/n487 ), .C(CLK), .Q(\U2/x[16][7] ), .QN(n97)
         );
  DF3 \U2/x_reg[15][0]  ( .D(\U2/n488 ), .C(CLK), .Q(\U2/x[15][0] ), .QN(n188)
         );
  DF3 \U2/x_reg[15][1]  ( .D(\U2/n489 ), .C(CLK), .Q(\U2/x[15][1] ), .QN(n187)
         );
  DF3 \U2/x_reg[15][2]  ( .D(\U2/n490 ), .C(CLK), .Q(\U2/x[15][2] ), .QN(n186)
         );
  DF3 \U2/x_reg[15][3]  ( .D(\U2/n491 ), .C(CLK), .Q(\U2/x[15][3] ), .QN(n185)
         );
  DF3 \U2/x_reg[15][4]  ( .D(\U2/n492 ), .C(CLK), .Q(\U2/x[15][4] ), .QN(n184)
         );
  DF3 \U2/x_reg[15][5]  ( .D(\U2/n493 ), .C(CLK), .Q(\U2/x[15][5] ), .QN(n183)
         );
  DF3 \U2/x_reg[15][6]  ( .D(\U2/n494 ), .C(CLK), .Q(\U2/x[15][6] ), .QN(n182)
         );
  DF3 \U2/x_reg[15][7]  ( .D(\U2/n495 ), .C(CLK), .Q(\U2/x[15][7] ), .QN(n181)
         );
  DF3 \U2/x_reg[14][0]  ( .D(\U2/n496 ), .C(CLK), .Q(\U2/x[14][0] ), .QN(n96)
         );
  DF3 \U2/x_reg[14][1]  ( .D(\U2/n497 ), .C(CLK), .Q(\U2/x[14][1] ), .QN(n95)
         );
  DF3 \U2/x_reg[14][2]  ( .D(\U2/n498 ), .C(CLK), .Q(\U2/x[14][2] ), .QN(n94)
         );
  DF3 \U2/x_reg[14][3]  ( .D(\U2/n499 ), .C(CLK), .Q(\U2/x[14][3] ), .QN(n93)
         );
  DF3 \U2/x_reg[14][4]  ( .D(\U2/n500 ), .C(CLK), .Q(\U2/x[14][4] ), .QN(n92)
         );
  DF3 \U2/x_reg[14][5]  ( .D(\U2/n501 ), .C(CLK), .Q(\U2/x[14][5] ), .QN(n91)
         );
  DF3 \U2/x_reg[14][6]  ( .D(\U2/n502 ), .C(CLK), .Q(\U2/x[14][6] ), .QN(n90)
         );
  DF3 \U2/x_reg[14][7]  ( .D(\U2/n503 ), .C(CLK), .Q(\U2/x[14][7] ), .QN(n89)
         );
  DF3 \U2/x_reg[13][0]  ( .D(\U2/n504 ), .C(CLK), .Q(\U2/x[13][0] ), .QN(n180)
         );
  DF3 \U2/x_reg[13][1]  ( .D(\U2/n505 ), .C(CLK), .Q(\U2/x[13][1] ), .QN(n153)
         );
  DF3 \U2/x_reg[13][2]  ( .D(\U2/n506 ), .C(CLK), .Q(\U2/x[13][2] ), .QN(n179)
         );
  DF3 \U2/x_reg[13][3]  ( .D(\U2/n507 ), .C(CLK), .Q(\U2/x[13][3] ), .QN(n178)
         );
  DF3 \U2/x_reg[13][4]  ( .D(\U2/n508 ), .C(CLK), .Q(\U2/x[13][4] ), .QN(n177)
         );
  DF3 \U2/x_reg[13][5]  ( .D(\U2/n509 ), .C(CLK), .Q(\U2/x[13][5] ), .QN(n176)
         );
  DF3 \U2/x_reg[13][6]  ( .D(\U2/n510 ), .C(CLK), .Q(\U2/x[13][6] ), .QN(n175)
         );
  DF3 \U2/x_reg[13][7]  ( .D(\U2/n511 ), .C(CLK), .Q(\U2/x[13][7] ), .QN(n174)
         );
  DF3 \U2/x_reg[12][0]  ( .D(\U2/n512 ), .C(CLK), .Q(\U2/x[12][0] ), .QN(n88)
         );
  DF3 \U2/x_reg[12][1]  ( .D(\U2/n513 ), .C(CLK), .Q(\U2/x[12][1] ), .QN(n59)
         );
  DF3 \U2/x_reg[12][2]  ( .D(\U2/n514 ), .C(CLK), .Q(\U2/x[12][2] ), .QN(n87)
         );
  DF3 \U2/x_reg[12][3]  ( .D(\U2/n515 ), .C(CLK), .Q(\U2/x[12][3] ), .QN(n86)
         );
  DF3 \U2/x_reg[12][4]  ( .D(\U2/n524 ), .C(CLK), .Q(\U2/x[12][4] ), .QN(n85)
         );
  DF3 \U2/x_reg[12][5]  ( .D(\U2/n525 ), .C(CLK), .Q(\U2/x[12][5] ), .QN(n84)
         );
  DF3 \U2/x_reg[12][6]  ( .D(\U2/n526 ), .C(CLK), .Q(\U2/x[12][6] ), .QN(n83)
         );
  DF3 \U2/x_reg[12][7]  ( .D(\U2/n527 ), .C(CLK), .Q(\U2/x[12][7] ), .QN(n82)
         );
  DF3 \U2/x_reg[11][0]  ( .D(\U2/n528 ), .C(CLK), .Q(\U2/x[11][0] ), .QN(n173)
         );
  DF3 \U2/x_reg[11][1]  ( .D(\U2/n529 ), .C(CLK), .Q(\U2/x[11][1] ), .QN(n152)
         );
  DF3 \U2/x_reg[11][2]  ( .D(\U2/n530 ), .C(CLK), .Q(\U2/x[11][2] ), .QN(n172)
         );
  DF3 \U2/x_reg[11][3]  ( .D(\U2/n531 ), .C(CLK), .Q(\U2/x[11][3] ), .QN(n171)
         );
  DF3 \U2/x_reg[11][4]  ( .D(\U2/n532 ), .C(CLK), .Q(\U2/x[11][4] ), .QN(n170)
         );
  DF3 \U2/x_reg[11][5]  ( .D(\U2/n533 ), .C(CLK), .Q(\U2/x[11][5] ), .QN(n169)
         );
  DF3 \U2/x_reg[11][6]  ( .D(\U2/n534 ), .C(CLK), .Q(\U2/x[11][6] ), .QN(n168)
         );
  DF3 \U2/x_reg[11][7]  ( .D(\U2/n535 ), .C(CLK), .Q(\U2/x[11][7] ), .QN(n167)
         );
  DF3 \U2/x_reg[10][0]  ( .D(\U2/n536 ), .C(CLK), .Q(\U2/x[10][0] ), .QN(n81)
         );
  DF3 \U2/x_reg[10][1]  ( .D(\U2/n537 ), .C(CLK), .Q(\U2/x[10][1] ), .QN(n58)
         );
  DF3 \U2/x_reg[10][2]  ( .D(\U2/n538 ), .C(CLK), .Q(\U2/x[10][2] ), .QN(n80)
         );
  DF3 \U2/x_reg[10][3]  ( .D(\U2/n539 ), .C(CLK), .Q(\U2/x[10][3] ), .QN(n79)
         );
  DF3 \U2/x_reg[10][4]  ( .D(\U2/n540 ), .C(CLK), .Q(\U2/x[10][4] ), .QN(n78)
         );
  DF3 \U2/x_reg[10][5]  ( .D(\U2/n541 ), .C(CLK), .Q(\U2/x[10][5] ), .QN(n77)
         );
  DF3 \U2/x_reg[10][6]  ( .D(\U2/n542 ), .C(CLK), .Q(\U2/x[10][6] ), .QN(n76)
         );
  DF3 \U2/x_reg[10][7]  ( .D(\U2/n543 ), .C(CLK), .Q(\U2/x[10][7] ), .QN(n75)
         );
  DF3 \U2/x_reg[9][0]  ( .D(\U2/n544 ), .C(CLK), .Q(\U2/x[9][0] ), .QN(n166)
         );
  DF3 \U2/x_reg[9][1]  ( .D(\U2/n545 ), .C(CLK), .Q(\U2/x[9][1] ), .QN(n151)
         );
  DF3 \U2/x_reg[9][2]  ( .D(\U2/n546 ), .C(CLK), .Q(\U2/x[9][2] ), .QN(n165)
         );
  DF3 \U2/x_reg[9][3]  ( .D(\U2/n547 ), .C(CLK), .Q(\U2/x[9][3] ), .QN(n164)
         );
  DF3 \U2/x_reg[9][4]  ( .D(\U2/n548 ), .C(CLK), .Q(\U2/x[9][4] ), .QN(n163)
         );
  DF3 \U2/x_reg[9][5]  ( .D(\U2/n549 ), .C(CLK), .Q(\U2/x[9][5] ), .QN(n162)
         );
  DF3 \U2/x_reg[9][6]  ( .D(\U2/n550 ), .C(CLK), .Q(\U2/x[9][6] ), .QN(n161)
         );
  DF3 \U2/x_reg[9][7]  ( .D(\U2/n551 ), .C(CLK), .Q(\U2/x[9][7] ), .QN(n160)
         );
  DF3 \U2/x_reg[8][0]  ( .D(\U2/n552 ), .C(CLK), .Q(\U2/x[8][0] ), .QN(n74) );
  DF3 \U2/x_reg[8][1]  ( .D(\U2/n553 ), .C(CLK), .Q(\U2/x[8][1] ), .QN(n57) );
  DF3 \U2/x_reg[8][2]  ( .D(\U2/n554 ), .C(CLK), .Q(\U2/x[8][2] ), .QN(n73) );
  DF3 \U2/x_reg[8][3]  ( .D(\U2/n555 ), .C(CLK), .Q(\U2/x[8][3] ), .QN(n72) );
  DF3 \U2/x_reg[8][4]  ( .D(\U2/n556 ), .C(CLK), .Q(\U2/x[8][4] ), .QN(n71) );
  DF3 \U2/x_reg[8][5]  ( .D(\U2/n557 ), .C(CLK), .Q(\U2/x[8][5] ), .QN(n70) );
  DF3 \U2/x_reg[8][6]  ( .D(\U2/n558 ), .C(CLK), .Q(\U2/x[8][6] ), .QN(n69) );
  DF3 \U2/x_reg[8][7]  ( .D(\U2/n559 ), .C(CLK), .Q(\U2/x[8][7] ), .QN(n68) );
  DF3 \U2/x_reg[7][0]  ( .D(\U2/n560 ), .C(CLK), .QN(n126) );
  DF3 \U2/x_reg[7][1]  ( .D(\U2/n561 ), .C(CLK), .QN(n122) );
  DF3 \U2/x_reg[7][2]  ( .D(\U2/n562 ), .C(CLK), .QN(n129) );
  DF3 \U2/x_reg[7][3]  ( .D(\U2/n563 ), .C(CLK), .QN(n132) );
  DF3 \U2/x_reg[7][4]  ( .D(\U2/n564 ), .C(CLK), .QN(n138) );
  DF3 \U2/x_reg[7][5]  ( .D(\U2/n565 ), .C(CLK), .QN(n135) );
  DF3 \U2/x_reg[7][6]  ( .D(\U2/n566 ), .C(CLK), .QN(n146) );
  DF3 \U2/x_reg[7][7]  ( .D(\U2/n567 ), .C(CLK), .QN(n142) );
  DF3 \U2/x_reg[6][0]  ( .D(\U2/n568 ), .C(CLK), .QN(n36) );
  DF3 \U2/x_reg[6][1]  ( .D(\U2/n569 ), .C(CLK), .QN(n33) );
  DF3 \U2/x_reg[6][2]  ( .D(\U2/n570 ), .C(CLK), .QN(n39) );
  DF3 \U2/x_reg[6][3]  ( .D(\U2/n571 ), .C(CLK), .QN(n43) );
  DF3 \U2/x_reg[6][4]  ( .D(\U2/n572 ), .C(CLK), .QN(n50) );
  DF3 \U2/x_reg[6][5]  ( .D(\U2/n573 ), .C(CLK), .QN(n47) );
  DF3 \U2/x_reg[6][6]  ( .D(\U2/n574 ), .C(CLK), .QN(n55) );
  DF3 \U2/x_reg[6][7]  ( .D(\U2/n575 ), .C(CLK), .QN(n53) );
  DF3 \U2/x_reg[5][0]  ( .D(\U2/n576 ), .C(CLK), .QN(n125) );
  DF3 \U2/x_reg[5][1]  ( .D(\U2/n577 ), .C(CLK), .QN(n123) );
  DF3 \U2/x_reg[5][2]  ( .D(\U2/n578 ), .C(CLK), .QN(n128) );
  DF3 \U2/x_reg[5][3]  ( .D(\U2/n579 ), .C(CLK), .QN(n131) );
  DF3 \U2/x_reg[5][4]  ( .D(\U2/n580 ), .C(CLK), .QN(n139) );
  DF3 \U2/x_reg[5][5]  ( .D(\U2/n581 ), .C(CLK), .QN(n136) );
  DF3 \U2/x_reg[5][6]  ( .D(\U2/n582 ), .C(CLK), .QN(n147) );
  DF3 \U2/x_reg[5][7]  ( .D(\U2/n583 ), .C(CLK), .QN(n143) );
  DF3 \U2/x_reg[4][0]  ( .D(\U2/n584 ), .C(CLK), .QN(n35) );
  DF3 \U2/x_reg[4][1]  ( .D(\U2/n585 ), .C(CLK), .QN(n34) );
  DF3 \U2/x_reg[4][2]  ( .D(\U2/n586 ), .C(CLK), .QN(n38) );
  DF3 \U2/x_reg[4][3]  ( .D(\U2/n587 ), .C(CLK), .QN(n42) );
  DF3 \U2/x_reg[4][4]  ( .D(\U2/n588 ), .C(CLK), .QN(n51) );
  DF3 \U2/x_reg[4][5]  ( .D(\U2/n589 ), .C(CLK), .QN(n48) );
  DF3 \U2/x_reg[4][6]  ( .D(\U2/n590 ), .C(CLK), .QN(n29) );
  DF3 \U2/x_reg[4][7]  ( .D(\U2/n591 ), .C(CLK), .QN(n27) );
  DF3 \U2/x_reg[3][0]  ( .D(\U2/n32 ), .C(CLK), .Q(\U2/x[3][0] ), .QN(n208) );
  DF3 \U2/x_reg[3][1]  ( .D(\U2/n31 ), .C(CLK), .Q(\U2/x[3][1] ), .QN(n207) );
  DF3 \U2/x_reg[3][2]  ( .D(\U2/n30 ), .C(CLK), .Q(\U2/x[3][2] ), .QN(n214) );
  DF3 \U2/x_reg[3][3]  ( .D(\U2/n29 ), .C(CLK), .Q(\U2/x[3][3] ), .QN(n213) );
  DF3 \U2/x_reg[3][4]  ( .D(\U2/n28 ), .C(CLK), .Q(\U2/x[3][4] ), .QN(n212) );
  DF3 \U2/x_reg[3][5]  ( .D(\U2/n27 ), .C(CLK), .Q(\U2/x[3][5] ), .QN(n211) );
  DF3 \U2/x_reg[3][6]  ( .D(\U2/n26 ), .C(CLK), .Q(\U2/x[3][6] ), .QN(n210) );
  DF3 \U2/x_reg[3][7]  ( .D(\U2/n25 ), .C(CLK), .Q(\U2/x[3][7] ), .QN(n209) );
  DF3 \U2/x_reg[2][0]  ( .D(\U2/n24 ), .C(CLK), .Q(\U2/x[2][0] ) );
  DF3 \U2/x_reg[2][1]  ( .D(\U2/n23 ), .C(CLK), .Q(\U2/x[2][1] ) );
  DF3 \U2/x_reg[2][2]  ( .D(\U2/n22 ), .C(CLK), .Q(\U2/x[2][2] ) );
  DF3 \U2/x_reg[2][3]  ( .D(\U2/n21 ), .C(CLK), .Q(\U2/x[2][3] ) );
  DF3 \U2/x_reg[2][4]  ( .D(\U2/n20 ), .C(CLK), .Q(\U2/x[2][4] ) );
  DF3 \U2/x_reg[2][5]  ( .D(\U2/n19 ), .C(CLK), .Q(\U2/x[2][5] ) );
  DF3 \U2/x_reg[2][6]  ( .D(\U2/n18 ), .C(CLK), .Q(\U2/x[2][6] ) );
  DF3 \U2/x_reg[2][7]  ( .D(\U2/n17 ), .C(CLK), .Q(\U2/x[2][7] ) );
  DF3 \U2/x_reg[1][0]  ( .D(\U2/n15 ), .C(CLK), .Q(\U2/x[1][0] ) );
  DF3 \U2/x_reg[1][1]  ( .D(\U2/n13 ), .C(CLK), .Q(\U2/x[1][1] ) );
  DF3 \U2/x_reg[1][2]  ( .D(\U2/n11 ), .C(CLK), .Q(\U2/x[1][2] ) );
  DF3 \U2/x_reg[1][3]  ( .D(\U2/n9 ), .C(CLK), .Q(\U2/x[1][3] ) );
  DF3 \U2/x_reg[1][4]  ( .D(\U2/n7 ), .C(CLK), .Q(\U2/x[1][4] ) );
  DF3 \U2/x_reg[1][5]  ( .D(\U2/n5 ), .C(CLK), .Q(\U2/x[1][5] ) );
  DF3 \U2/x_reg[1][6]  ( .D(\U2/n3 ), .C(CLK), .Q(\U2/x[1][6] ) );
  DF3 \U2/x_reg[1][7]  ( .D(\U2/n1 ), .C(CLK), .Q(\U2/x[1][7] ) );
  DF3 \U2/x_reg[0][0]  ( .D(\U2/n16 ), .C(CLK), .Q(\U2/x[0][0] ) );
  DF3 \U2/x_reg[0][1]  ( .D(\U2/n14 ), .C(CLK), .Q(\U2/x[0][1] ) );
  DF3 \U2/x_reg[0][2]  ( .D(\U2/n12 ), .C(CLK), .Q(\U2/x[0][2] ) );
  DF3 \U2/x_reg[0][3]  ( .D(\U2/n10 ), .C(CLK), .Q(\U2/x[0][3] ) );
  DF3 \U2/x_reg[0][4]  ( .D(\U2/n8 ), .C(CLK), .Q(\U2/x[0][4] ) );
  DF3 \U2/x_reg[0][5]  ( .D(\U2/n6 ), .C(CLK), .Q(\U2/x[0][5] ) );
  DF3 \U2/x_reg[0][6]  ( .D(\U2/n4 ), .C(CLK), .Q(\U2/x[0][6] ) );
  DF3 \U2/x_reg[0][7]  ( .D(\U2/n2 ), .C(CLK), .Q(\U2/x[0][7] ) );
  DF3 \U4/ACCU_reg[19]  ( .D(\U4/N46 ), .C(CLK), .Q(Accu_out[19]) );
  DF3 \U4/ACCU_reg[18]  ( .D(\U4/N45 ), .C(CLK), .Q(Accu_out[18]) );
  DF3 \U4/ACCU_reg[17]  ( .D(\U4/N44 ), .C(CLK), .Q(Accu_out[17]) );
  DF3 \U4/ACCU_reg[16]  ( .D(\U4/N43 ), .C(CLK), .Q(Accu_out[16]) );
  DF3 \U4/ACCU_reg[15]  ( .D(\U4/N42 ), .C(CLK), .Q(Accu_out[15]) );
  DF3 \U4/ACCU_reg[14]  ( .D(\U4/N41 ), .C(CLK), .Q(Accu_out[14]) );
  DF3 \U4/ACCU_reg[13]  ( .D(\U4/N40 ), .C(CLK), .Q(Accu_out[13]), .QN(n8) );
  DF3 \U4/ACCU_reg[12]  ( .D(\U4/N39 ), .C(CLK), .Q(Accu_out[12]) );
  DF3 \U4/ACCU_reg[11]  ( .D(\U4/N38 ), .C(CLK), .Q(\U4/Accu_out[11] ) );
  DF3 \U4/ACCU_reg[10]  ( .D(\U4/N37 ), .C(CLK), .Q(\U4/Accu_out[10] ) );
  DF3 \U4/ACCU_reg[9]  ( .D(\U4/N36 ), .C(CLK), .Q(\U4/Accu_out[9] ) );
  DF3 \U4/ACCU_reg[8]  ( .D(\U4/N35 ), .C(CLK), .Q(\U4/Accu_out[8] ) );
  DF3 \U4/ACCU_reg[7]  ( .D(\U4/N34 ), .C(CLK), .Q(\U4/Accu_out[7] ) );
  DF3 \U4/ACCU_reg[6]  ( .D(\U4/N33 ), .C(CLK), .Q(\U4/Accu_out[6] ) );
  DF3 \U4/ACCU_reg[5]  ( .D(\U4/N32 ), .C(CLK), .Q(\U4/Accu_out[5] ) );
  DF3 \U4/ACCU_reg[4]  ( .D(\U4/N31 ), .C(CLK), .Q(\U4/Accu_out[4] ) );
  DF3 \U4/ACCU_reg[3]  ( .D(\U4/N30 ), .C(CLK), .Q(\U4/Accu_out[3] ) );
  DF3 \U4/ACCU_reg[2]  ( .D(\U4/N29 ), .C(CLK), .Q(\U4/Accu_out[2] ) );
  DF3 \U4/ACCU_reg[1]  ( .D(\U4/N28 ), .C(CLK), .Q(\U4/Accu_out[1] ) );
  DF3 \U4/ACCU_reg[0]  ( .D(\U4/N27 ), .C(CLK), .Q(\U4/Accu_out[0] ) );
  OAI212 \U5/U17  ( .A(\U5/n19 ), .B(\U5/n1 ), .C(\U5/n10 ), .Q(\U5/n20 ) );
  OAI212 \U5/U15  ( .A(\U5/n18 ), .B(\U5/n1 ), .C(\U5/n9 ), .Q(\U5/n21 ) );
  OAI212 \U5/U13  ( .A(\U5/n17 ), .B(\U5/n1 ), .C(\U5/n8 ), .Q(\U5/n22 ) );
  OAI212 \U5/U11  ( .A(\U5/n16 ), .B(\U5/n1 ), .C(\U5/n7 ), .Q(\U5/n23 ) );
  OAI212 \U5/U9  ( .A(\U5/n15 ), .B(\U5/n1 ), .C(\U5/n6 ), .Q(\U5/n24 ) );
  OAI212 \U5/U7  ( .A(\U5/n14 ), .B(\U5/n1 ), .C(\U5/n5 ), .Q(\U5/n25 ) );
  OAI212 \U5/U5  ( .A(\U5/n13 ), .B(\U5/n1 ), .C(\U5/n4 ), .Q(\U5/n26 ) );
  OAI212 \U5/U3  ( .A(\U5/n12 ), .B(\U5/n1 ), .C(\U5/n2 ), .Q(\U5/n27 ) );
  DF3 \U5/Buff_out_reg[0]  ( .D(\U5/n27 ), .C(CLK), .Q(Filter_Out[0]), .QN(
        \U5/n12 ) );
  DF3 \U5/Buff_out_reg[1]  ( .D(\U5/n26 ), .C(CLK), .Q(Filter_Out[1]), .QN(
        \U5/n13 ) );
  DF3 \U5/Buff_out_reg[2]  ( .D(\U5/n25 ), .C(CLK), .Q(Filter_Out[2]), .QN(
        \U5/n14 ) );
  DF3 \U5/Buff_out_reg[3]  ( .D(\U5/n24 ), .C(CLK), .Q(Filter_Out[3]), .QN(
        \U5/n15 ) );
  DF3 \U5/Buff_out_reg[4]  ( .D(\U5/n23 ), .C(CLK), .Q(Filter_Out[4]), .QN(
        \U5/n16 ) );
  DF3 \U5/Buff_out_reg[5]  ( .D(\U5/n22 ), .C(CLK), .Q(Filter_Out[5]), .QN(
        \U5/n17 ) );
  DF3 \U5/Buff_out_reg[6]  ( .D(\U5/n21 ), .C(CLK), .Q(Filter_Out[6]), .QN(
        \U5/n18 ) );
  DF3 \U5/Buff_out_reg[7]  ( .D(\U5/n20 ), .C(CLK), .Q(Filter_Out[7]), .QN(
        \U5/n19 ) );
  OAI212 \U6/U13  ( .A(\U6/n33 ), .B(n121), .C(n233), .Q(\U6/n36 ) );
  OAI212 \U6/U6  ( .A(\U6/n13 ), .B(\U1/n7 ), .C(\U6/n29 ), .Q(\U6/n42 ) );
  DFC3 \U6/cpt_current_reg[3]  ( .D(\U6/n40 ), .C(CLK), .RN(n263), .Q(\U6/n47 ), .QN(n31) );
  DFC3 \U6/cpt_current_reg[2]  ( .D(\U6/n39 ), .C(CLK), .RN(n263), .QN(n19) );
  DFC3 \U6/cpt_current_reg[1]  ( .D(\U6/n38 ), .C(CLK), .RN(n263), .Q(n223), 
        .QN(\U6/n33 ) );
  DFC3 \U6/cpt_current_reg[4]  ( .D(\U6/n42 ), .C(CLK), .RN(n263), .Q(\U6/n48 ) );
  DFC3 \U6/current_state_reg[2]  ( .D(\U6/n41 ), .C(CLK), .RN(n263), .Q(n149), 
        .QN(\U6/n14 ) );
  DFC3 \U6/current_state_reg[1]  ( .D(\U6/n7 ), .C(CLK), .RN(n263), .Q(
        \U6/n50 ), .QN(n30) );
  DFC3 \U6/cpt_current_reg[0]  ( .D(\U6/n37 ), .C(CLK), .RN(n263), .Q(\U6/n4 ), 
        .QN(n121) );
  DFC3 \U6/current_state_reg[0]  ( .D(\U6/n10 ), .C(CLK), .RN(n263), .Q(
        \U6/n2 ) );
  OAI212 \U7/U10  ( .A(n56), .B(n148), .C(\U7/n12 ), .Q(ADC_Convstb) );
  OAI222 \U7/U4  ( .A(\U7/n2 ), .B(ack_F2ADC), .C(req_ADC2F), .D(\U7/n11 ), 
        .Q(\U7/n10 ) );
  DFC3 \U7/current_state_reg[1]  ( .D(\U7/n14 ), .C(CLK), .RN(n263), .Q(
        \U7/n2 ), .QN(n148) );
  DFC3 \U7/current_state_reg[2]  ( .D(\U7/n13 ), .C(CLK), .RN(n263), .Q(n56)
         );
  DFC3 \U7/current_state_reg[0]  ( .D(\U7/n15 ), .C(CLK), .RN(n263), .Q(n150), 
        .QN(\U7/n9 ) );
  DF3 \U8/current_state_reg  ( .D(\U8/N5 ), .C(CLK), .Q(\U8/current_state ), 
        .QN(DAC_WRb) );
  DF3 \U8/pre_req_F2DAC_reg  ( .D(\U8/n1 ), .C(CLK), .Q(\U8/pre_req_F2DAC ) );
  OAI212 \U9/U17  ( .A(\U9/n1 ), .B(\U9/n19 ), .C(\U9/n10 ), .Q(\U9/n20 ) );
  OAI212 \U9/U15  ( .A(\U9/n1 ), .B(\U9/n18 ), .C(\U9/n9 ), .Q(\U9/n21 ) );
  OAI212 \U9/U13  ( .A(\U9/n1 ), .B(\U9/n17 ), .C(\U9/n8 ), .Q(\U9/n22 ) );
  OAI212 \U9/U11  ( .A(\U9/n1 ), .B(\U9/n16 ), .C(\U9/n7 ), .Q(\U9/n23 ) );
  OAI212 \U9/U9  ( .A(\U9/n1 ), .B(\U9/n15 ), .C(\U9/n6 ), .Q(\U9/n24 ) );
  OAI212 \U9/U7  ( .A(\U9/n1 ), .B(\U9/n14 ), .C(\U9/n5 ), .Q(\U9/n25 ) );
  OAI212 \U9/U5  ( .A(\U9/n1 ), .B(\U9/n13 ), .C(\U9/n4 ), .Q(\U9/n26 ) );
  OAI212 \U9/U3  ( .A(\U9/n1 ), .B(\U9/n12 ), .C(\U9/n2 ), .Q(\U9/n27 ) );
  DF3 \U9/reg_reg[0]  ( .D(\U9/n27 ), .C(CLK), .Q(Filter_In_mem[0]), .QN(
        \U9/n12 ) );
  DF3 \U9/reg_reg[1]  ( .D(\U9/n26 ), .C(CLK), .Q(Filter_In_mem[1]), .QN(
        \U9/n13 ) );
  DF3 \U9/reg_reg[2]  ( .D(\U9/n25 ), .C(CLK), .Q(Filter_In_mem[2]), .QN(
        \U9/n14 ) );
  DF3 \U9/reg_reg[3]  ( .D(\U9/n24 ), .C(CLK), .Q(Filter_In_mem[3]), .QN(
        \U9/n15 ) );
  DF3 \U9/reg_reg[4]  ( .D(\U9/n23 ), .C(CLK), .Q(Filter_In_mem[4]), .QN(
        \U9/n16 ) );
  DF3 \U9/reg_reg[5]  ( .D(\U9/n22 ), .C(CLK), .Q(Filter_In_mem[5]), .QN(
        \U9/n17 ) );
  DF3 \U9/reg_reg[6]  ( .D(\U9/n21 ), .C(CLK), .Q(Filter_In_mem[6]), .QN(
        \U9/n18 ) );
  DF3 \U9/reg_reg[7]  ( .D(\U9/n20 ), .C(CLK), .Q(Filter_In_mem[7]), .QN(
        \U9/n19 ) );
  ADD32 \U3/mult_19/S3_2_6  ( .A(\U3/mult_19/ab[2][6] ), .B(
        \U3/mult_19/CARRYB[1][6] ), .CI(\U3/mult_19/ab[1][7] ), .CO(
        \U3/mult_19/CARRYB[2][6] ), .S(\U3/mult_19/SUMB[2][6] ) );
  ADD32 \U3/mult_19/S2_2_5  ( .A(\U3/mult_19/ab[2][5] ), .B(
        \U3/mult_19/CARRYB[1][5] ), .CI(\U3/mult_19/SUMB[1][6] ), .CO(
        \U3/mult_19/CARRYB[2][5] ), .S(\U3/mult_19/SUMB[2][5] ) );
  ADD32 \U3/mult_19/S2_2_4  ( .A(\U3/mult_19/ab[2][4] ), .B(
        \U3/mult_19/CARRYB[1][4] ), .CI(\U3/mult_19/SUMB[1][5] ), .CO(
        \U3/mult_19/CARRYB[2][4] ), .S(\U3/mult_19/SUMB[2][4] ) );
  ADD32 \U3/mult_19/S2_2_3  ( .A(\U3/mult_19/ab[2][3] ), .B(
        \U3/mult_19/CARRYB[1][3] ), .CI(\U3/mult_19/SUMB[1][4] ), .CO(
        \U3/mult_19/CARRYB[2][3] ), .S(\U3/mult_19/SUMB[2][3] ) );
  ADD32 \U3/mult_19/S2_2_2  ( .A(\U3/mult_19/ab[2][2] ), .B(
        \U3/mult_19/CARRYB[1][2] ), .CI(\U3/mult_19/SUMB[1][3] ), .CO(
        \U3/mult_19/CARRYB[2][2] ), .S(\U3/mult_19/SUMB[2][2] ) );
  ADD32 \U3/mult_19/S2_2_1  ( .A(\U3/mult_19/ab[2][1] ), .B(
        \U3/mult_19/CARRYB[1][1] ), .CI(\U3/mult_19/SUMB[1][2] ), .CO(
        \U3/mult_19/CARRYB[2][1] ), .S(\U3/mult_19/SUMB[2][1] ) );
  ADD32 \U3/mult_19/S1_2_0  ( .A(\U3/mult_19/ab[2][0] ), .B(
        \U3/mult_19/CARRYB[1][0] ), .CI(\U3/mult_19/SUMB[1][1] ), .CO(
        \U3/mult_19/CARRYB[2][0] ), .S(Mult_out[2]) );
  ADD32 \U3/mult_19/S3_3_6  ( .A(\U3/mult_19/ab[3][6] ), .B(
        \U3/mult_19/CARRYB[2][6] ), .CI(\U3/mult_19/ab[2][7] ), .CO(
        \U3/mult_19/CARRYB[3][6] ), .S(\U3/mult_19/SUMB[3][6] ) );
  ADD32 \U3/mult_19/S2_3_5  ( .A(\U3/mult_19/ab[3][5] ), .B(
        \U3/mult_19/CARRYB[2][5] ), .CI(\U3/mult_19/SUMB[2][6] ), .CO(
        \U3/mult_19/CARRYB[3][5] ), .S(\U3/mult_19/SUMB[3][5] ) );
  ADD32 \U3/mult_19/S2_3_4  ( .A(\U3/mult_19/ab[3][4] ), .B(
        \U3/mult_19/CARRYB[2][4] ), .CI(\U3/mult_19/SUMB[2][5] ), .CO(
        \U3/mult_19/CARRYB[3][4] ), .S(\U3/mult_19/SUMB[3][4] ) );
  ADD32 \U3/mult_19/S2_3_3  ( .A(\U3/mult_19/ab[3][3] ), .B(
        \U3/mult_19/CARRYB[2][3] ), .CI(\U3/mult_19/SUMB[2][4] ), .CO(
        \U3/mult_19/CARRYB[3][3] ), .S(\U3/mult_19/SUMB[3][3] ) );
  ADD32 \U3/mult_19/S2_3_2  ( .A(\U3/mult_19/ab[3][2] ), .B(
        \U3/mult_19/CARRYB[2][2] ), .CI(\U3/mult_19/SUMB[2][3] ), .CO(
        \U3/mult_19/CARRYB[3][2] ), .S(\U3/mult_19/SUMB[3][2] ) );
  ADD32 \U3/mult_19/S2_3_1  ( .A(\U3/mult_19/ab[3][1] ), .B(
        \U3/mult_19/CARRYB[2][1] ), .CI(\U3/mult_19/SUMB[2][2] ), .CO(
        \U3/mult_19/CARRYB[3][1] ), .S(\U3/mult_19/SUMB[3][1] ) );
  ADD32 \U3/mult_19/S1_3_0  ( .A(\U3/mult_19/ab[3][0] ), .B(
        \U3/mult_19/CARRYB[2][0] ), .CI(\U3/mult_19/SUMB[2][1] ), .CO(
        \U3/mult_19/CARRYB[3][0] ), .S(Mult_out[3]) );
  ADD32 \U3/mult_19/S3_4_6  ( .A(\U3/mult_19/ab[4][6] ), .B(
        \U3/mult_19/CARRYB[3][6] ), .CI(\U3/mult_19/ab[3][7] ), .CO(
        \U3/mult_19/CARRYB[4][6] ), .S(\U3/mult_19/SUMB[4][6] ) );
  ADD32 \U3/mult_19/S2_4_5  ( .A(\U3/mult_19/ab[4][5] ), .B(
        \U3/mult_19/CARRYB[3][5] ), .CI(\U3/mult_19/SUMB[3][6] ), .CO(
        \U3/mult_19/CARRYB[4][5] ), .S(\U3/mult_19/SUMB[4][5] ) );
  ADD32 \U3/mult_19/S2_4_4  ( .A(\U3/mult_19/ab[4][4] ), .B(
        \U3/mult_19/CARRYB[3][4] ), .CI(\U3/mult_19/SUMB[3][5] ), .CO(
        \U3/mult_19/CARRYB[4][4] ), .S(\U3/mult_19/SUMB[4][4] ) );
  ADD32 \U3/mult_19/S2_4_3  ( .A(\U3/mult_19/ab[4][3] ), .B(
        \U3/mult_19/CARRYB[3][3] ), .CI(\U3/mult_19/SUMB[3][4] ), .CO(
        \U3/mult_19/CARRYB[4][3] ), .S(\U3/mult_19/SUMB[4][3] ) );
  ADD32 \U3/mult_19/S2_4_2  ( .A(\U3/mult_19/ab[4][2] ), .B(
        \U3/mult_19/CARRYB[3][2] ), .CI(\U3/mult_19/SUMB[3][3] ), .CO(
        \U3/mult_19/CARRYB[4][2] ), .S(\U3/mult_19/SUMB[4][2] ) );
  ADD32 \U3/mult_19/S2_4_1  ( .A(\U3/mult_19/ab[4][1] ), .B(
        \U3/mult_19/CARRYB[3][1] ), .CI(\U3/mult_19/SUMB[3][2] ), .CO(
        \U3/mult_19/CARRYB[4][1] ), .S(\U3/mult_19/SUMB[4][1] ) );
  ADD32 \U3/mult_19/S1_4_0  ( .A(\U3/mult_19/ab[4][0] ), .B(
        \U3/mult_19/CARRYB[3][0] ), .CI(\U3/mult_19/SUMB[3][1] ), .CO(
        \U3/mult_19/CARRYB[4][0] ), .S(Mult_out[4]) );
  ADD32 \U3/mult_19/S3_5_6  ( .A(\U3/mult_19/ab[5][6] ), .B(
        \U3/mult_19/CARRYB[4][6] ), .CI(\U3/mult_19/ab[4][7] ), .CO(
        \U3/mult_19/CARRYB[5][6] ), .S(\U3/mult_19/SUMB[5][6] ) );
  ADD32 \U3/mult_19/S2_5_5  ( .A(\U3/mult_19/ab[5][5] ), .B(
        \U3/mult_19/CARRYB[4][5] ), .CI(\U3/mult_19/SUMB[4][6] ), .CO(
        \U3/mult_19/CARRYB[5][5] ), .S(\U3/mult_19/SUMB[5][5] ) );
  ADD32 \U3/mult_19/S2_5_4  ( .A(\U3/mult_19/ab[5][4] ), .B(
        \U3/mult_19/CARRYB[4][4] ), .CI(\U3/mult_19/SUMB[4][5] ), .CO(
        \U3/mult_19/CARRYB[5][4] ), .S(\U3/mult_19/SUMB[5][4] ) );
  ADD32 \U3/mult_19/S2_5_3  ( .A(\U3/mult_19/ab[5][3] ), .B(
        \U3/mult_19/CARRYB[4][3] ), .CI(\U3/mult_19/SUMB[4][4] ), .CO(
        \U3/mult_19/CARRYB[5][3] ), .S(\U3/mult_19/SUMB[5][3] ) );
  ADD32 \U3/mult_19/S2_5_2  ( .A(\U3/mult_19/ab[5][2] ), .B(
        \U3/mult_19/CARRYB[4][2] ), .CI(\U3/mult_19/SUMB[4][3] ), .CO(
        \U3/mult_19/CARRYB[5][2] ), .S(\U3/mult_19/SUMB[5][2] ) );
  ADD32 \U3/mult_19/S2_5_1  ( .A(\U3/mult_19/ab[5][1] ), .B(
        \U3/mult_19/CARRYB[4][1] ), .CI(\U3/mult_19/SUMB[4][2] ), .CO(
        \U3/mult_19/CARRYB[5][1] ), .S(\U3/mult_19/SUMB[5][1] ) );
  ADD32 \U3/mult_19/S1_5_0  ( .A(\U3/mult_19/ab[5][0] ), .B(
        \U3/mult_19/CARRYB[4][0] ), .CI(\U3/mult_19/SUMB[4][1] ), .CO(
        \U3/mult_19/CARRYB[5][0] ), .S(Mult_out[5]) );
  ADD32 \U3/mult_19/S3_6_6  ( .A(\U3/mult_19/ab[6][6] ), .B(
        \U3/mult_19/CARRYB[5][6] ), .CI(\U3/mult_19/ab[5][7] ), .CO(
        \U3/mult_19/CARRYB[6][6] ), .S(\U3/mult_19/SUMB[6][6] ) );
  ADD32 \U3/mult_19/S2_6_5  ( .A(\U3/mult_19/ab[6][5] ), .B(
        \U3/mult_19/CARRYB[5][5] ), .CI(\U3/mult_19/SUMB[5][6] ), .CO(
        \U3/mult_19/CARRYB[6][5] ), .S(\U3/mult_19/SUMB[6][5] ) );
  ADD32 \U3/mult_19/S2_6_4  ( .A(\U3/mult_19/ab[6][4] ), .B(
        \U3/mult_19/CARRYB[5][4] ), .CI(\U3/mult_19/SUMB[5][5] ), .CO(
        \U3/mult_19/CARRYB[6][4] ), .S(\U3/mult_19/SUMB[6][4] ) );
  ADD32 \U3/mult_19/S2_6_3  ( .A(\U3/mult_19/ab[6][3] ), .B(
        \U3/mult_19/CARRYB[5][3] ), .CI(\U3/mult_19/SUMB[5][4] ), .CO(
        \U3/mult_19/CARRYB[6][3] ), .S(\U3/mult_19/SUMB[6][3] ) );
  ADD32 \U3/mult_19/S2_6_2  ( .A(\U3/mult_19/ab[6][2] ), .B(
        \U3/mult_19/CARRYB[5][2] ), .CI(\U3/mult_19/SUMB[5][3] ), .CO(
        \U3/mult_19/CARRYB[6][2] ), .S(\U3/mult_19/SUMB[6][2] ) );
  ADD32 \U3/mult_19/S2_6_1  ( .A(\U3/mult_19/ab[6][1] ), .B(
        \U3/mult_19/CARRYB[5][1] ), .CI(\U3/mult_19/SUMB[5][2] ), .CO(
        \U3/mult_19/CARRYB[6][1] ), .S(\U3/mult_19/SUMB[6][1] ) );
  ADD32 \U3/mult_19/S1_6_0  ( .A(\U3/mult_19/ab[6][0] ), .B(
        \U3/mult_19/CARRYB[5][0] ), .CI(\U3/mult_19/SUMB[5][1] ), .CO(
        \U3/mult_19/CARRYB[6][0] ), .S(Mult_out[6]) );
  ADD32 \U3/mult_19/S5_6  ( .A(\U3/mult_19/ab[7][6] ), .B(
        \U3/mult_19/CARRYB[6][6] ), .CI(\U3/mult_19/ab[6][7] ), .CO(
        \U3/mult_19/CARRYB[7][6] ), .S(\U3/mult_19/SUMB[7][6] ) );
  ADD32 \U3/mult_19/S4_5  ( .A(\U3/mult_19/ab[7][5] ), .B(
        \U3/mult_19/CARRYB[6][5] ), .CI(\U3/mult_19/SUMB[6][6] ), .CO(
        \U3/mult_19/CARRYB[7][5] ), .S(\U3/mult_19/SUMB[7][5] ) );
  ADD32 \U3/mult_19/S4_4  ( .A(\U3/mult_19/ab[7][4] ), .B(
        \U3/mult_19/CARRYB[6][4] ), .CI(\U3/mult_19/SUMB[6][5] ), .CO(
        \U3/mult_19/CARRYB[7][4] ), .S(\U3/mult_19/SUMB[7][4] ) );
  ADD32 \U3/mult_19/S4_3  ( .A(\U3/mult_19/ab[7][3] ), .B(
        \U3/mult_19/CARRYB[6][3] ), .CI(\U3/mult_19/SUMB[6][4] ), .CO(
        \U3/mult_19/CARRYB[7][3] ), .S(\U3/mult_19/SUMB[7][3] ) );
  ADD32 \U3/mult_19/S4_2  ( .A(\U3/mult_19/ab[7][2] ), .B(
        \U3/mult_19/CARRYB[6][2] ), .CI(\U3/mult_19/SUMB[6][3] ), .CO(
        \U3/mult_19/CARRYB[7][2] ), .S(\U3/mult_19/SUMB[7][2] ) );
  ADD32 \U3/mult_19/S4_1  ( .A(\U3/mult_19/ab[7][1] ), .B(
        \U3/mult_19/CARRYB[6][1] ), .CI(\U3/mult_19/SUMB[6][2] ), .CO(
        \U3/mult_19/CARRYB[7][1] ), .S(\U3/mult_19/SUMB[7][1] ) );
  ADD32 \U3/mult_19/S4_0  ( .A(\U3/mult_19/ab[7][0] ), .B(
        \U3/mult_19/CARRYB[6][0] ), .CI(\U3/mult_19/SUMB[6][1] ), .CO(
        \U3/mult_19/CARRYB[7][0] ), .S(Mult_out[7]) );
  ADD32 \U4/add_27_aco/U1_1  ( .A(\U4/N49 ), .B(Mult_out[1]), .CI(
        \U4/add_27_aco/carry [1]), .CO(\U4/add_27_aco/carry [2]), .S(\U4/N7 )
         );
  ADD32 \U4/add_27_aco/U1_2  ( .A(\U4/N50 ), .B(Mult_out[2]), .CI(
        \U4/add_27_aco/carry [2]), .CO(\U4/add_27_aco/carry [3]), .S(\U4/N8 )
         );
  ADD32 \U4/add_27_aco/U1_3  ( .A(\U4/N51 ), .B(Mult_out[3]), .CI(
        \U4/add_27_aco/carry [3]), .CO(\U4/add_27_aco/carry [4]), .S(\U4/N9 )
         );
  ADD32 \U4/add_27_aco/U1_4  ( .A(\U4/N52 ), .B(Mult_out[4]), .CI(
        \U4/add_27_aco/carry [4]), .CO(\U4/add_27_aco/carry [5]), .S(\U4/N10 )
         );
  ADD32 \U4/add_27_aco/U1_5  ( .A(\U4/N53 ), .B(Mult_out[5]), .CI(
        \U4/add_27_aco/carry [5]), .CO(\U4/add_27_aco/carry [6]), .S(\U4/N11 )
         );
  ADD32 \U4/add_27_aco/U1_6  ( .A(\U4/N54 ), .B(Mult_out[6]), .CI(
        \U4/add_27_aco/carry [6]), .CO(\U4/add_27_aco/carry [7]), .S(\U4/N12 )
         );
  ADD32 \U4/add_27_aco/U1_7  ( .A(\U4/N55 ), .B(Mult_out[7]), .CI(
        \U4/add_27_aco/carry [7]), .CO(\U4/add_27_aco/carry [8]), .S(\U4/N13 )
         );
  ADD32 \U4/add_27_aco/U1_8  ( .A(\U4/N56 ), .B(Mult_out[8]), .CI(
        \U4/add_27_aco/carry [8]), .CO(\U4/add_27_aco/carry [9]), .S(\U4/N14 )
         );
  ADD32 \U4/add_27_aco/U1_9  ( .A(\U4/N57 ), .B(Mult_out[9]), .CI(
        \U4/add_27_aco/carry [9]), .CO(\U4/add_27_aco/carry [10]), .S(\U4/N15 ) );
  ADD32 \U4/add_27_aco/U1_10  ( .A(\U4/N58 ), .B(Mult_out[10]), .CI(
        \U4/add_27_aco/carry [10]), .CO(\U4/add_27_aco/carry [11]), .S(
        \U4/N16 ) );
  ADD32 \U4/add_27_aco/U1_11  ( .A(\U4/N59 ), .B(Mult_out[11]), .CI(
        \U4/add_27_aco/carry [11]), .CO(\U4/add_27_aco/carry [12]), .S(
        \U4/N17 ) );
  ADD32 \U4/add_27_aco/U1_12  ( .A(\U4/N60 ), .B(Mult_out[12]), .CI(
        \U4/add_27_aco/carry [12]), .CO(\U4/add_27_aco/carry [13]), .S(
        \U4/N18 ) );
  ADD32 \U4/add_27_aco/U1_13  ( .A(\U4/N61 ), .B(Mult_out[13]), .CI(
        \U4/add_27_aco/carry [13]), .CO(\U4/add_27_aco/carry [14]), .S(
        \U4/N19 ) );
  ADD32 \U4/add_27_aco/U1_14  ( .A(\U4/N62 ), .B(Mult_out[14]), .CI(
        \U4/add_27_aco/carry [14]), .CO(\U4/add_27_aco/carry [15]), .S(
        \U4/N20 ) );
  ADD32 \U4/add_27_aco/U1_15  ( .A(\U4/N63 ), .B(Mult_out[15]), .CI(
        \U4/add_27_aco/carry [15]), .CO(\U4/add_27_aco/carry [16]), .S(
        \U4/N21 ) );
  OAI212 \U3/mult_19/FS_1/U37  ( .A(\U3/mult_19/FS_1/n12 ), .B(
        \U3/mult_19/FS_1/n31 ), .C(\U3/mult_19/FS_1/n13 ), .Q(
        \U3/mult_19/FS_1/n9 ) );
  XOR31 \U3/mult_19/FS_1/U28  ( .A(\U3/mult_19/A2[11] ), .B(
        \U3/mult_19/A1[11] ), .C(\U3/mult_19/FS_1/n28 ), .Q(Mult_out[13]) );
  OAI212 \U3/mult_19/FS_1/U27  ( .A(\U3/mult_19/FS_1/n13 ), .B(
        \U3/mult_19/FS_1/n22 ), .C(\U3/mult_19/FS_1/n11 ), .Q(
        \U3/mult_19/FS_1/n27 ) );
  OAI212 \U3/mult_19/FS_1/U26  ( .A(\U3/mult_19/FS_1/n23 ), .B(
        \U3/mult_19/FS_1/n37 ), .C(\U3/mult_19/FS_1/n26 ), .Q(
        \U3/mult_19/FS_1/n20 ) );
  OAI212 \U3/mult_19/FS_1/U25  ( .A(\U3/mult_19/A1[11] ), .B(
        \U3/mult_19/FS_1/n20 ), .C(\U3/mult_19/A2[11] ), .Q(
        \U3/mult_19/FS_1/n25 ) );
  XOR31 \U3/mult_19/FS_1/U21  ( .A(\U3/mult_19/A2[12] ), .B(
        \U3/mult_19/A1[12] ), .C(\U3/mult_19/FS_1/n33 ), .Q(Mult_out[14]) );
  OAI212 \U3/mult_19/FS_1/U20  ( .A(\U3/mult_19/A1[12] ), .B(
        \U3/mult_19/FS_1/n33 ), .C(\U3/mult_19/A2[12] ), .Q(
        \U3/mult_19/FS_1/n18 ) );
  OAI212 \U3/mult_19/FS_1/U15  ( .A(\U3/mult_19/FS_1/n12 ), .B(
        \U3/mult_19/FS_1/n13 ), .C(\U3/mult_19/FS_1/n14 ), .Q(Mult_out[10]) );
  NOR22 U12 ( .A(\U6/n44 ), .B(\U6/n33 ), .Q(n229) );
  NAND22 U13 ( .A(\U3/mult_19/ab[0][2] ), .B(\U3/mult_19/ab[1][1] ), .Q(n3) );
  INV3 U14 ( .A(n3), .Q(\U3/mult_19/CARRYB[1][1] ) );
  MUX22 U15 ( .A(\U2/n523 ), .B(\U2/n522 ), .S(\U6/n29 ), .Q(\U3/mult_19/n64 )
         );
  NAND22 U16 ( .A(\U3/mult_19/CARRYB[7][3] ), .B(\U3/mult_19/SUMB[7][4] ), .Q(
        n4) );
  INV3 U17 ( .A(n4), .Q(\U3/mult_19/A2[10] ) );
  NOR30 U18 ( .A(n149), .B(\U6/n2 ), .C(n30), .Q(Buff_OE) );
  MUX22 U19 ( .A(\U2/n613 ), .B(\U2/n612 ), .S(\U6/n29 ), .Q(\U3/mult_19/n65 )
         );
  NAND22 U20 ( .A(\U3/mult_19/CARRYB[7][4] ), .B(\U3/mult_19/SUMB[7][5] ), .Q(
        n5) );
  INV3 U21 ( .A(n5), .Q(\U3/mult_19/A2[11] ) );
  NOR20 U22 ( .A(\U6/n16 ), .B(\U6/n2 ), .Q(Delay_Line_sample_shift) );
  XNR21 U23 ( .A(n11), .B(\U3/mult_19/A1[7] ), .Q(Mult_out[9]) );
  NAND22 U24 ( .A(\U3/mult_19/ab[0][7] ), .B(\U3/mult_19/ab[1][6] ), .Q(n6) );
  INV3 U25 ( .A(n6), .Q(\U3/mult_19/CARRYB[1][6] ) );
  XNR31 U26 ( .A(\U3/mult_19/FS_1/n29 ), .B(\U3/mult_19/A2[10] ), .C(
        \U3/mult_19/A1[10] ), .Q(Mult_out[12]) );
  NAND22 U27 ( .A(\U3/mult_19/CARRYB[7][1] ), .B(\U3/mult_19/SUMB[7][2] ), .Q(
        n7) );
  INV3 U28 ( .A(n7), .Q(\U3/mult_19/A2[8] ) );
  MUX22 U29 ( .A(\U2/n701 ), .B(\U2/n700 ), .S(\U6/n29 ), .Q(\U3/mult_19/n83 )
         );
  AOI211 U30 ( .A(\U6/n2 ), .B(ack_F2ADC), .C(n8), .Q(\U4/N61 ) );
  MUX22 U31 ( .A(\U2/n351 ), .B(\U2/n350 ), .S(\U6/n29 ), .Q(\U3/mult_19/n62 )
         );
  NAND22 U32 ( .A(\U3/mult_19/ab[0][1] ), .B(\U3/mult_19/ab[1][0] ), .Q(n9) );
  INV3 U33 ( .A(n9), .Q(\U3/mult_19/CARRYB[1][0] ) );
  XOR21 U34 ( .A(\U3/mult_19/FS_1/n17 ), .B(n13), .Q(Mult_out[15]) );
  NAND22 U35 ( .A(\U3/mult_19/ab[0][6] ), .B(\U3/mult_19/ab[1][5] ), .Q(n10)
         );
  INV3 U36 ( .A(n10), .Q(\U3/mult_19/CARRYB[1][5] ) );
  AOI311 U37 ( .A(n56), .B(\U7/n9 ), .C(n148), .D(RESET), .Q(\U9/n11 ) );
  NAND22 U38 ( .A(\U3/mult_19/CARRYB[7][0] ), .B(\U3/mult_19/SUMB[7][1] ), .Q(
        n11) );
  INV3 U39 ( .A(n11), .Q(\U3/mult_19/A2[7] ) );
  OAI212 U40 ( .A(\U3/mult_19/A2[9] ), .B(\U3/mult_19/A1[9] ), .C(
        \U3/mult_19/FS_1/n11 ), .Q(\U3/mult_19/FS_1/n10 ) );
  NAND22 U41 ( .A(\U3/mult_19/CARRYB[7][5] ), .B(\U3/mult_19/SUMB[7][6] ), .Q(
        n12) );
  INV3 U42 ( .A(n12), .Q(\U3/mult_19/A2[12] ) );
  NOR31 U43 ( .A(\U4/add_27_aco/n18 ), .B(\U4/mult_add_27_aco/PROD_not[16] ), 
        .C(\U4/mult_add_27_aco/PROD_not[17] ), .Q(\U4/add_27_aco/carry [18])
         );
  IMUX21 U44 ( .A(\U1/n51 ), .B(\U1/n18 ), .S(Rom_Address[2]), .Q(\U1/n48 ) );
  IMAJ31 U45 ( .A(\U3/mult_19/FS_1/n9 ), .B(\U3/mult_19/A2[9] ), .C(
        \U3/mult_19/A1[9] ), .Q(\U3/mult_19/FS_1/n29 ) );
  NAND22 U46 ( .A(\U3/mult_19/CARRYB[7][6] ), .B(\U3/mult_19/ab[7][7] ), .Q(
        n13) );
  AOI211 U47 ( .A(\U6/n31 ), .B(req_ADC2F), .C(Delay_Line_sample_shift), .Q(
        n14) );
  INV3 U48 ( .A(n14), .Q(\U6/n41 ) );
  XOR21 U49 ( .A(\U4/mult_add_27_aco/PROD_not[0] ), .B(Mult_out[0]), .Q(n228)
         );
  NOR21 U50 ( .A(RESET), .B(n228), .Q(\U4/N27 ) );
  NOR21 U51 ( .A(RESET), .B(n225), .Q(\U4/N43 ) );
  NOR21 U52 ( .A(RESET), .B(n226), .Q(\U4/N44 ) );
  NOR21 U53 ( .A(RESET), .B(n227), .Q(\U4/N45 ) );
  NOR21 U54 ( .A(n232), .B(n231), .Q(\U2/n716 ) );
  NAND22 U55 ( .A(\U2/n716 ), .B(\U2/n717 ), .Q(\U2/n357 ) );
  NAND22 U56 ( .A(\U2/n716 ), .B(\U2/n720 ), .Q(\U2/n358 ) );
  CLKIN3 U57 ( .A(n230), .Q(\U1/n12 ) );
  INV3 U58 ( .A(n229), .Q(\U2/n280 ) );
  INV3 U59 ( .A(\U2/n723 ), .Q(\U2/n269 ) );
  BUF2 U60 ( .A(Rom_Address[0]), .Q(n230) );
  XOR21 U61 ( .A(\U4/mult_add_27_aco/PROD_not[19] ), .B(
        \U4/add_27_aco/carry [19]), .Q(n224) );
  NAND22 U62 ( .A(\U3/mult_19/A2[8] ), .B(\U3/mult_19/A1[8] ), .Q(
        \U3/mult_19/FS_1/n13 ) );
  NAND20 U63 ( .A(\U2/n718 ), .B(\U2/n724 ), .Q(\U2/n726 ) );
  INV1 U64 ( .A(\U3/mult_19/ab[1][2] ), .Q(\U3/mult_19/n70 ) );
  INV2 U65 ( .A(\U3/mult_19/ab[0][4] ), .Q(\U3/mult_19/n79 ) );
  NAND22 U66 ( .A(\U2/n716 ), .B(\U2/n719 ), .Q(\U2/n359 ) );
  INV3 U67 ( .A(\U2/n734 ), .Q(\U2/n276 ) );
  CLKIN1 U68 ( .A(n231), .Q(\U2/n278 ) );
  INV3 U69 ( .A(\U4/add_27_aco/carry [16]), .Q(\U4/add_27_aco/n18 ) );
  OAI222 U70 ( .A(n15), .B(\U2/n358 ), .C(n32), .D(\U2/n359 ), .Q(\U2/n682 )
         );
  INV3 U71 ( .A(Delay_Line_out[1]), .Q(\U3/mult_19/n75 ) );
  AOI221 U72 ( .A(\U2/n272 ), .B(\U2/x[12][1] ), .C(\U2/n273 ), .D(
        \U2/x[13][1] ), .Q(\U2/n697 ) );
  AOI221 U73 ( .A(\U2/n274 ), .B(\U2/x[10][1] ), .C(\U2/n275 ), .D(
        \U2/x[11][1] ), .Q(\U2/n698 ) );
  AOI221 U74 ( .A(\U2/n276 ), .B(\U2/x[8][1] ), .C(\U2/n277 ), .D(\U2/x[9][1] ), .Q(\U2/n699 ) );
  NOR20 U75 ( .A(n121), .B(\U6/n44 ), .Q(Rom_Address[0]) );
  OAI211 U76 ( .A(\U3/mult_19/FS_1/n23 ), .B(\U3/mult_19/FS_1/n29 ), .C(
        \U3/mult_19/FS_1/n26 ), .Q(\U3/mult_19/FS_1/n28 ) );
  NOR20 U77 ( .A(\U3/mult_19/A1[8] ), .B(\U3/mult_19/A2[8] ), .Q(
        \U3/mult_19/FS_1/n31 ) );
  NOR20 U78 ( .A(\U3/mult_19/A1[8] ), .B(\U3/mult_19/FS_1/n39 ), .Q(
        \U3/mult_19/FS_1/n16 ) );
  INV1 U79 ( .A(\U3/mult_19/FS_1/n12 ), .Q(\U3/mult_19/FS_1/n39 ) );
  OAI220 U80 ( .A(\U3/mult_19/A1[11] ), .B(\U3/mult_19/A2[11] ), .C(
        \U3/mult_19/A1[8] ), .D(\U3/mult_19/A2[8] ), .Q(\U3/mult_19/FS_1/n24 )
         );
  NAND20 U81 ( .A(\U2/n717 ), .B(\U2/n724 ), .Q(\U2/n727 ) );
  CLKIN3 U82 ( .A(\U2/n741 ), .Q(\U2/n270 ) );
  NAND21 U83 ( .A(\U2/n738 ), .B(\U2/n717 ), .Q(\U2/n741 ) );
  CLKIN3 U84 ( .A(\U2/n725 ), .Q(\U2/n268 ) );
  NAND20 U85 ( .A(\U2/n724 ), .B(\U2/n719 ), .Q(\U2/n725 ) );
  NAND20 U86 ( .A(\U2/n720 ), .B(\U2/n724 ), .Q(\U2/n723 ) );
  CLKIN3 U87 ( .A(\U2/n737 ), .Q(\U2/n273 ) );
  NAND21 U88 ( .A(\U2/n738 ), .B(\U2/n720 ), .Q(\U2/n737 ) );
  NOR20 U89 ( .A(\U3/mult_19/n88 ), .B(\U3/mult_19/n75 ), .Q(
        \U3/mult_19/ab[1][3] ) );
  NOR20 U90 ( .A(\U3/mult_19/n90 ), .B(\U3/mult_19/n75 ), .Q(
        \U3/mult_19/ab[1][1] ) );
  NOR20 U91 ( .A(\U3/mult_19/n91 ), .B(\U3/mult_19/n75 ), .Q(
        \U3/mult_19/ab[1][0] ) );
  NOR20 U92 ( .A(\U3/mult_19/n89 ), .B(\U3/mult_19/n75 ), .Q(
        \U3/mult_19/ab[1][2] ) );
  NOR20 U93 ( .A(\U3/mult_19/n89 ), .B(\U3/mult_19/n83 ), .Q(
        \U3/mult_19/ab[0][2] ) );
  NOR20 U94 ( .A(\U3/mult_19/n90 ), .B(\U3/mult_19/n83 ), .Q(
        \U3/mult_19/ab[0][1] ) );
  NOR20 U95 ( .A(\U3/mult_19/n88 ), .B(\U3/mult_19/n83 ), .Q(
        \U3/mult_19/ab[0][3] ) );
  NOR20 U96 ( .A(\U3/mult_19/n87 ), .B(\U3/mult_19/n83 ), .Q(
        \U3/mult_19/ab[0][4] ) );
  NOR20 U97 ( .A(\U3/mult_19/n84 ), .B(\U3/mult_19/n75 ), .Q(
        \U3/mult_19/ab[1][7] ) );
  INV2 U98 ( .A(n231), .Q(\U1/n7 ) );
  NAND21 U99 ( .A(Rom_Address[4]), .B(n231), .Q(\U1/n20 ) );
  NOR20 U100 ( .A(\U1/n40 ), .B(n231), .Q(\U1/n28 ) );
  NAND30 U101 ( .A(Rom_Address[4]), .B(\U2/n280 ), .C(n230), .Q(\U1/n26 ) );
  AOI220 U102 ( .A(\U1/n23 ), .B(\U1/n7 ), .C(\U1/n24 ), .D(n230), .Q(\U1/n22 ) );
  OAI210 U103 ( .A(n231), .B(Rom_Address[4]), .C(\U1/n20 ), .Q(\U1/n37 ) );
  NAND20 U104 ( .A(n230), .B(n233), .Q(\U1/n30 ) );
  OAI210 U105 ( .A(n230), .B(\U1/n25 ), .C(\U1/n26 ), .Q(\U1/n23 ) );
  NOR20 U106 ( .A(\U3/mult_19/n91 ), .B(\U3/mult_19/n83 ), .Q(Mult_out[0]) );
  AOI210 U107 ( .A(n230), .B(\U2/n280 ), .C(\U1/n20 ), .Q(\U1/n43 ) );
  OAI310 U108 ( .A(\U2/n280 ), .B(n231), .C(\U1/n2 ), .D(\U1/n26 ), .Q(
        \U1/n50 ) );
  NAND20 U109 ( .A(\U2/n733 ), .B(\U2/n719 ), .Q(\U2/n734 ) );
  OAI221 U110 ( .A(n125), .B(\U2/n358 ), .C(n35), .D(\U2/n359 ), .Q(\U2/n714 )
         );
  OAI221 U111 ( .A(n127), .B(\U2/n358 ), .C(n37), .D(\U2/n359 ), .Q(\U2/n704 )
         );
  OAI220 U112 ( .A(n130), .B(\U2/n358 ), .C(n40), .D(\U2/n359 ), .Q(\U2/n660 )
         );
  OAI220 U113 ( .A(n128), .B(\U2/n358 ), .C(n38), .D(\U2/n359 ), .Q(\U2/n670 )
         );
  OAI221 U114 ( .A(n126), .B(\U2/n356 ), .C(n36), .D(n235), .Q(\U2/n715 ) );
  OAI221 U115 ( .A(n21), .B(\U2/n356 ), .C(n16), .D(n235), .Q(\U2/n705 ) );
  OAI221 U116 ( .A(n20), .B(\U2/n356 ), .C(n124), .D(n235), .Q(\U2/n683 ) );
  OAI220 U117 ( .A(n22), .B(\U2/n356 ), .C(n41), .D(n235), .Q(\U2/n661 ) );
  OAI220 U118 ( .A(n129), .B(\U2/n356 ), .C(n39), .D(n235), .Q(\U2/n671 ) );
  XNR20 U119 ( .A(\U4/N65 ), .B(\U4/add_27_aco/carry [17]), .Q(n226) );
  XNR20 U120 ( .A(\U4/N66 ), .B(\U4/add_27_aco/carry [18]), .Q(n227) );
  OAI211 U121 ( .A(n229), .B(\U1/n12 ), .C(\U1/n29 ), .Q(\U1/n32 ) );
  NAND21 U122 ( .A(n229), .B(\U1/n12 ), .Q(\U1/n29 ) );
  NAND20 U123 ( .A(n229), .B(n230), .Q(\U1/n40 ) );
  OAI220 U124 ( .A(n133), .B(\U2/n358 ), .C(n44), .D(\U2/n359 ), .Q(\U2/n638 )
         );
  OAI220 U125 ( .A(n131), .B(\U2/n358 ), .C(n42), .D(\U2/n359 ), .Q(\U2/n648 )
         );
  OAI220 U126 ( .A(n23), .B(\U2/n356 ), .C(n45), .D(n235), .Q(\U2/n639 ) );
  OAI220 U127 ( .A(n132), .B(\U2/n356 ), .C(n43), .D(n235), .Q(\U2/n649 ) );
  XNR20 U128 ( .A(\U4/N64 ), .B(\U4/add_27_aco/carry [16]), .Q(n225) );
  OAI210 U129 ( .A(n229), .B(\U1/n7 ), .C(\U1/n29 ), .Q(\U1/n51 ) );
  AOI220 U130 ( .A(\U2/n270 ), .B(\U2/x[14][1] ), .C(\U2/n271 ), .D(
        \U2/x[15][1] ), .Q(\U2/n696 ) );
  AOI220 U131 ( .A(\U2/n274 ), .B(\U2/x[10][0] ), .C(\U2/n275 ), .D(
        \U2/x[11][0] ), .Q(\U2/n730 ) );
  AOI220 U132 ( .A(\U2/n276 ), .B(\U2/x[8][0] ), .C(\U2/n277 ), .D(
        \U2/x[9][0] ), .Q(\U2/n731 ) );
  AOI220 U133 ( .A(\U2/n270 ), .B(\U2/x[14][0] ), .C(\U2/n271 ), .D(
        \U2/x[15][0] ), .Q(\U2/n728 ) );
  AOI220 U134 ( .A(\U2/n274 ), .B(\U2/x[26][2] ), .C(\U2/n275 ), .D(
        \U2/x[27][2] ), .Q(\U2/n666 ) );
  AOI220 U135 ( .A(\U2/n276 ), .B(\U2/x[24][2] ), .C(\U2/n277 ), .D(
        \U2/x[25][2] ), .Q(\U2/n667 ) );
  AOI220 U136 ( .A(\U2/n270 ), .B(\U2/x[30][2] ), .C(\U2/n271 ), .D(
        \U2/x[31][2] ), .Q(\U2/n664 ) );
  AOI220 U137 ( .A(\U2/n276 ), .B(\U2/x[8][2] ), .C(\U2/n277 ), .D(
        \U2/x[9][2] ), .Q(\U2/n677 ) );
  AOI220 U138 ( .A(\U2/n274 ), .B(\U2/x[10][2] ), .C(\U2/n275 ), .D(
        \U2/x[11][2] ), .Q(\U2/n676 ) );
  AOI220 U139 ( .A(\U2/n270 ), .B(\U2/x[14][2] ), .C(\U2/n271 ), .D(
        \U2/x[15][2] ), .Q(\U2/n674 ) );
  AOI220 U140 ( .A(\U2/n274 ), .B(\U2/x[26][3] ), .C(\U2/n275 ), .D(
        \U2/x[27][3] ), .Q(\U2/n644 ) );
  AOI220 U141 ( .A(\U2/n276 ), .B(\U2/x[24][3] ), .C(\U2/n277 ), .D(
        \U2/x[25][3] ), .Q(\U2/n645 ) );
  AOI220 U142 ( .A(\U2/n270 ), .B(\U2/x[30][3] ), .C(\U2/n271 ), .D(
        \U2/x[31][3] ), .Q(\U2/n642 ) );
  AOI220 U143 ( .A(\U2/n274 ), .B(\U2/x[10][3] ), .C(\U2/n275 ), .D(
        \U2/x[11][3] ), .Q(\U2/n654 ) );
  AOI220 U144 ( .A(\U2/n276 ), .B(\U2/x[8][3] ), .C(\U2/n277 ), .D(
        \U2/x[9][3] ), .Q(\U2/n655 ) );
  AOI220 U145 ( .A(\U2/n270 ), .B(\U2/x[14][3] ), .C(\U2/n271 ), .D(
        \U2/x[15][3] ), .Q(\U2/n652 ) );
  AOI220 U146 ( .A(\U2/n272 ), .B(\U2/x[12][0] ), .C(\U2/n273 ), .D(
        \U2/x[13][0] ), .Q(\U2/n729 ) );
  AOI220 U147 ( .A(\U2/n272 ), .B(\U2/x[28][2] ), .C(\U2/n273 ), .D(
        \U2/x[29][2] ), .Q(\U2/n665 ) );
  AOI220 U148 ( .A(\U2/n272 ), .B(\U2/x[12][2] ), .C(\U2/n273 ), .D(
        \U2/x[13][2] ), .Q(\U2/n675 ) );
  AOI220 U149 ( .A(\U2/n272 ), .B(\U2/x[28][3] ), .C(\U2/n273 ), .D(
        \U2/x[29][3] ), .Q(\U2/n643 ) );
  AOI220 U150 ( .A(\U2/n272 ), .B(\U2/x[12][3] ), .C(\U2/n273 ), .D(
        \U2/x[13][3] ), .Q(\U2/n653 ) );
  XOR20 U151 ( .A(\U3/mult_19/SUMB[7][1] ), .B(\U3/mult_19/CARRYB[7][0] ), .Q(
        Mult_out[8]) );
  AOI220 U152 ( .A(\U2/n268 ), .B(\U2/x[0][1] ), .C(\U2/n269 ), .D(
        \U2/x[1][1] ), .Q(\U2/n695 ) );
  AOI220 U153 ( .A(\U2/n268 ), .B(\U2/x[0][0] ), .C(\U2/n269 ), .D(
        \U2/x[1][0] ), .Q(\U2/n722 ) );
  AOI220 U154 ( .A(\U2/n266 ), .B(\U2/x[18][2] ), .C(\U2/n267 ), .D(
        \U2/x[19][2] ), .Q(\U2/n662 ) );
  AOI220 U155 ( .A(\U2/n268 ), .B(\U2/x[16][2] ), .C(\U2/n269 ), .D(
        \U2/x[17][2] ), .Q(\U2/n663 ) );
  AOI220 U156 ( .A(\U2/n268 ), .B(\U2/x[0][2] ), .C(\U2/n269 ), .D(
        \U2/x[1][2] ), .Q(\U2/n673 ) );
  AOI220 U157 ( .A(\U2/n266 ), .B(\U2/x[2][2] ), .C(\U2/n267 ), .D(
        \U2/x[3][2] ), .Q(\U2/n672 ) );
  AOI220 U158 ( .A(\U2/n266 ), .B(\U2/x[18][3] ), .C(\U2/n267 ), .D(
        \U2/x[19][3] ), .Q(\U2/n640 ) );
  AOI220 U159 ( .A(\U2/n268 ), .B(\U2/x[16][3] ), .C(\U2/n269 ), .D(
        \U2/x[17][3] ), .Q(\U2/n641 ) );
  AOI220 U160 ( .A(\U2/n274 ), .B(\U2/x[26][4] ), .C(\U2/n275 ), .D(
        \U2/x[27][4] ), .Q(\U2/n622 ) );
  AOI220 U161 ( .A(\U2/n276 ), .B(\U2/x[24][4] ), .C(\U2/n277 ), .D(
        \U2/x[25][4] ), .Q(\U2/n623 ) );
  AOI220 U162 ( .A(\U2/n270 ), .B(\U2/x[30][4] ), .C(\U2/n271 ), .D(
        \U2/x[31][4] ), .Q(\U2/n620 ) );
  AOI220 U163 ( .A(\U2/n274 ), .B(\U2/x[10][4] ), .C(\U2/n275 ), .D(
        \U2/x[11][4] ), .Q(\U2/n632 ) );
  AOI220 U164 ( .A(\U2/n276 ), .B(\U2/x[8][4] ), .C(\U2/n277 ), .D(
        \U2/x[9][4] ), .Q(\U2/n633 ) );
  AOI220 U165 ( .A(\U2/n270 ), .B(\U2/x[14][4] ), .C(\U2/n271 ), .D(
        \U2/x[15][4] ), .Q(\U2/n630 ) );
  AOI220 U166 ( .A(\U2/n274 ), .B(\U2/x[26][5] ), .C(\U2/n275 ), .D(
        \U2/x[27][5] ), .Q(\U2/n600 ) );
  AOI220 U167 ( .A(\U2/n276 ), .B(\U2/x[24][5] ), .C(\U2/n277 ), .D(
        \U2/x[25][5] ), .Q(\U2/n601 ) );
  AOI220 U168 ( .A(\U2/n270 ), .B(\U2/x[30][5] ), .C(\U2/n271 ), .D(
        \U2/x[31][5] ), .Q(\U2/n598 ) );
  AOI220 U169 ( .A(\U2/n274 ), .B(\U2/x[10][5] ), .C(\U2/n275 ), .D(
        \U2/x[11][5] ), .Q(\U2/n610 ) );
  AOI220 U170 ( .A(\U2/n276 ), .B(\U2/x[8][5] ), .C(\U2/n277 ), .D(
        \U2/x[9][5] ), .Q(\U2/n611 ) );
  AOI220 U171 ( .A(\U2/n270 ), .B(\U2/x[14][5] ), .C(\U2/n271 ), .D(
        \U2/x[15][5] ), .Q(\U2/n608 ) );
  AOI220 U172 ( .A(\U2/n266 ), .B(\U2/x[18][5] ), .C(\U2/n267 ), .D(
        \U2/x[19][5] ), .Q(\U2/n596 ) );
  AOI220 U173 ( .A(\U2/n268 ), .B(\U2/x[16][5] ), .C(\U2/n269 ), .D(
        \U2/x[17][5] ), .Q(\U2/n597 ) );
  AOI220 U174 ( .A(\U2/n272 ), .B(\U2/x[28][4] ), .C(\U2/n273 ), .D(
        \U2/x[29][4] ), .Q(\U2/n621 ) );
  AOI220 U175 ( .A(\U2/n272 ), .B(\U2/x[12][4] ), .C(\U2/n273 ), .D(
        \U2/x[13][4] ), .Q(\U2/n631 ) );
  AOI220 U176 ( .A(\U2/n272 ), .B(\U2/x[28][5] ), .C(\U2/n273 ), .D(
        \U2/x[29][5] ), .Q(\U2/n599 ) );
  AOI220 U177 ( .A(\U2/n272 ), .B(\U2/x[12][5] ), .C(\U2/n273 ), .D(
        \U2/x[13][5] ), .Q(\U2/n609 ) );
  AOI220 U178 ( .A(\U2/n266 ), .B(\U2/x[2][3] ), .C(\U2/n267 ), .D(
        \U2/x[3][3] ), .Q(\U2/n650 ) );
  AOI220 U179 ( .A(\U2/n268 ), .B(\U2/x[0][3] ), .C(\U2/n269 ), .D(
        \U2/x[1][3] ), .Q(\U2/n651 ) );
  AOI220 U180 ( .A(\U2/n266 ), .B(\U2/x[18][4] ), .C(\U2/n267 ), .D(
        \U2/x[19][4] ), .Q(\U2/n618 ) );
  AOI220 U181 ( .A(\U2/n268 ), .B(\U2/x[16][4] ), .C(\U2/n269 ), .D(
        \U2/x[17][4] ), .Q(\U2/n619 ) );
  AOI220 U182 ( .A(\U2/n266 ), .B(\U2/x[2][4] ), .C(\U2/n267 ), .D(
        \U2/x[3][4] ), .Q(\U2/n628 ) );
  AOI220 U183 ( .A(\U2/n268 ), .B(\U2/x[0][4] ), .C(\U2/n269 ), .D(
        \U2/x[1][4] ), .Q(\U2/n629 ) );
  AOI220 U184 ( .A(\U2/n266 ), .B(\U2/x[2][5] ), .C(\U2/n267 ), .D(
        \U2/x[3][5] ), .Q(\U2/n606 ) );
  AOI220 U185 ( .A(\U2/n268 ), .B(\U2/x[0][5] ), .C(\U2/n269 ), .D(
        \U2/x[1][5] ), .Q(\U2/n607 ) );
  AOI220 U186 ( .A(\U2/n266 ), .B(\U2/x[18][6] ), .C(\U2/n267 ), .D(
        \U2/x[19][6] ), .Q(\U2/n382 ) );
  AOI220 U187 ( .A(\U2/n268 ), .B(\U2/x[16][6] ), .C(\U2/n269 ), .D(
        \U2/x[17][6] ), .Q(\U2/n383 ) );
  AOI220 U188 ( .A(\U2/n266 ), .B(\U2/x[2][6] ), .C(\U2/n267 ), .D(
        \U2/x[3][6] ), .Q(\U2/n516 ) );
  AOI220 U189 ( .A(\U2/n268 ), .B(\U2/x[0][6] ), .C(\U2/n269 ), .D(
        \U2/x[1][6] ), .Q(\U2/n517 ) );
  AOI220 U190 ( .A(\U2/n274 ), .B(\U2/x[26][6] ), .C(\U2/n275 ), .D(
        \U2/x[27][6] ), .Q(\U2/n386 ) );
  AOI220 U191 ( .A(\U2/n276 ), .B(\U2/x[24][6] ), .C(\U2/n277 ), .D(
        \U2/x[25][6] ), .Q(\U2/n387 ) );
  AOI220 U192 ( .A(\U2/n270 ), .B(\U2/x[30][6] ), .C(\U2/n271 ), .D(
        \U2/x[31][6] ), .Q(\U2/n384 ) );
  AOI220 U193 ( .A(\U2/n274 ), .B(\U2/x[10][6] ), .C(\U2/n275 ), .D(
        \U2/x[11][6] ), .Q(\U2/n520 ) );
  AOI220 U194 ( .A(\U2/n276 ), .B(\U2/x[8][6] ), .C(\U2/n277 ), .D(
        \U2/x[9][6] ), .Q(\U2/n521 ) );
  AOI220 U195 ( .A(\U2/n270 ), .B(\U2/x[14][6] ), .C(\U2/n271 ), .D(
        \U2/x[15][6] ), .Q(\U2/n518 ) );
  AOI220 U196 ( .A(\U2/n274 ), .B(\U2/x[26][7] ), .C(\U2/n275 ), .D(
        \U2/x[27][7] ), .Q(\U2/n364 ) );
  AOI220 U197 ( .A(\U2/n276 ), .B(\U2/x[24][7] ), .C(\U2/n277 ), .D(
        \U2/x[25][7] ), .Q(\U2/n365 ) );
  AOI220 U198 ( .A(\U2/n270 ), .B(\U2/x[30][7] ), .C(\U2/n271 ), .D(
        \U2/x[31][7] ), .Q(\U2/n362 ) );
  AOI220 U199 ( .A(\U2/n272 ), .B(\U2/x[28][6] ), .C(\U2/n273 ), .D(
        \U2/x[29][6] ), .Q(\U2/n385 ) );
  AOI220 U200 ( .A(\U2/n272 ), .B(\U2/x[12][6] ), .C(\U2/n273 ), .D(
        \U2/x[13][6] ), .Q(\U2/n519 ) );
  AOI220 U201 ( .A(\U2/n266 ), .B(\U2/x[18][7] ), .C(\U2/n267 ), .D(
        \U2/x[19][7] ), .Q(\U2/n360 ) );
  AOI220 U202 ( .A(\U2/n268 ), .B(\U2/x[16][7] ), .C(\U2/n269 ), .D(
        \U2/x[17][7] ), .Q(\U2/n361 ) );
  AOI220 U203 ( .A(\U2/n268 ), .B(\U2/x[0][7] ), .C(\U2/n269 ), .D(
        \U2/x[1][7] ), .Q(\U2/n371 ) );
  AOI220 U204 ( .A(\U2/n266 ), .B(\U2/x[2][7] ), .C(\U2/n267 ), .D(
        \U2/x[3][7] ), .Q(\U2/n370 ) );
  AOI220 U205 ( .A(\U2/n276 ), .B(\U2/x[8][7] ), .C(\U2/n277 ), .D(
        \U2/x[9][7] ), .Q(\U2/n375 ) );
  AOI220 U206 ( .A(\U2/n274 ), .B(\U2/x[10][7] ), .C(\U2/n275 ), .D(
        \U2/x[11][7] ), .Q(\U2/n374 ) );
  AOI220 U207 ( .A(\U2/n270 ), .B(\U2/x[14][7] ), .C(\U2/n271 ), .D(
        \U2/x[15][7] ), .Q(\U2/n372 ) );
  AOI220 U208 ( .A(\U2/n272 ), .B(\U2/x[28][7] ), .C(\U2/n273 ), .D(
        \U2/x[29][7] ), .Q(\U2/n363 ) );
  AOI220 U209 ( .A(\U2/n272 ), .B(\U2/x[12][7] ), .C(\U2/n273 ), .D(
        \U2/x[13][7] ), .Q(\U2/n373 ) );
  NAND20 U210 ( .A(n229), .B(n121), .Q(\U6/n43 ) );
  NAND30 U211 ( .A(\U6/n4 ), .B(n19), .C(n229), .Q(\U6/n35 ) );
  NAND30 U212 ( .A(\U6/n2 ), .B(\U6/n14 ), .C(\U6/n50 ), .Q(\U6/n23 ) );
  OAI210 U213 ( .A(\U6/n50 ), .B(\U6/n2 ), .C(\U6/n23 ), .Q(\U6/n31 ) );
  NAND33 U214 ( .A(\U6/n14 ), .B(n30), .C(\U6/n2 ), .Q(\U6/n44 ) );
  INV3 U215 ( .A(\U3/mult_19/FS_1/n27 ), .Q(\U3/mult_19/FS_1/n37 ) );
  INV3 U216 ( .A(n250), .Q(n260) );
  INV3 U217 ( .A(n249), .Q(n259) );
  INV3 U218 ( .A(n249), .Q(n258) );
  INV3 U219 ( .A(n249), .Q(n257) );
  INV3 U220 ( .A(n250), .Q(n256) );
  INV3 U221 ( .A(\U2/n286 ), .Q(n255) );
  INV3 U222 ( .A(n249), .Q(n254) );
  INV3 U223 ( .A(n250), .Q(n253) );
  INV3 U224 ( .A(n250), .Q(n252) );
  INV3 U225 ( .A(n249), .Q(n251) );
  INV3 U226 ( .A(Rom_out[7]), .Q(\U3/mult_19/n84 ) );
  NAND22 U227 ( .A(\U3/mult_19/A2[7] ), .B(\U3/mult_19/A1[7] ), .Q(
        \U3/mult_19/FS_1/n12 ) );
  AOI211 U228 ( .A(\U3/mult_19/FS_1/n33 ), .B(\U3/mult_19/A1[12] ), .C(
        \U3/mult_19/FS_1/n32 ), .Q(\U3/mult_19/FS_1/n17 ) );
  INV3 U229 ( .A(\U3/mult_19/FS_1/n18 ), .Q(\U3/mult_19/FS_1/n32 ) );
  BUF2 U230 ( .A(\U2/n357 ), .Q(n235) );
  IMUX21 U231 ( .A(\U3/mult_19/FS_1/n15 ), .B(\U3/mult_19/FS_1/n16 ), .S(
        \U3/mult_19/A2[8] ), .Q(\U3/mult_19/FS_1/n14 ) );
  XNR21 U232 ( .A(\U3/mult_19/A1[8] ), .B(\U3/mult_19/FS_1/n12 ), .Q(
        \U3/mult_19/FS_1/n15 ) );
  INV3 U233 ( .A(\U3/mult_19/FS_1/n19 ), .Q(\U3/mult_19/FS_1/n33 ) );
  AOI2111 U234 ( .A(\U3/mult_19/FS_1/n20 ), .B(\U3/mult_19/A1[11] ), .C(
        \U3/mult_19/FS_1/n34 ), .D(\U3/mult_19/FS_1/n21 ), .Q(
        \U3/mult_19/FS_1/n19 ) );
  NOR40 U235 ( .A(\U3/mult_19/FS_1/n22 ), .B(\U3/mult_19/FS_1/n12 ), .C(
        \U3/mult_19/FS_1/n23 ), .D(\U3/mult_19/FS_1/n24 ), .Q(
        \U3/mult_19/FS_1/n21 ) );
  INV3 U236 ( .A(\U3/mult_19/FS_1/n25 ), .Q(\U3/mult_19/FS_1/n34 ) );
  NOR21 U237 ( .A(\U3/mult_19/A2[10] ), .B(\U3/mult_19/A1[10] ), .Q(
        \U3/mult_19/FS_1/n23 ) );
  NAND22 U238 ( .A(\U3/mult_19/A2[9] ), .B(\U3/mult_19/A1[9] ), .Q(
        \U3/mult_19/FS_1/n11 ) );
  NOR21 U239 ( .A(\U3/mult_19/A2[9] ), .B(\U3/mult_19/A1[9] ), .Q(
        \U3/mult_19/FS_1/n22 ) );
  NAND22 U240 ( .A(\U3/mult_19/A2[10] ), .B(\U3/mult_19/A1[10] ), .Q(
        \U3/mult_19/FS_1/n26 ) );
  INV3 U241 ( .A(\U1/n16 ), .Q(\U1/n6 ) );
  INV3 U242 ( .A(n248), .Q(n244) );
  INV3 U243 ( .A(n245), .Q(n243) );
  INV3 U244 ( .A(n246), .Q(n242) );
  INV3 U245 ( .A(n246), .Q(n241) );
  INV3 U246 ( .A(n245), .Q(n240) );
  INV3 U247 ( .A(n245), .Q(n239) );
  INV3 U248 ( .A(n248), .Q(n238) );
  INV3 U249 ( .A(n246), .Q(n237) );
  BUF2 U250 ( .A(n250), .Q(n261) );
  BUF2 U251 ( .A(n249), .Q(n262) );
  XOR21 U252 ( .A(\U3/mult_19/SUMB[7][3] ), .B(\U3/mult_19/CARRYB[7][2] ), .Q(
        \U3/mult_19/A1[8] ) );
  XOR21 U253 ( .A(\U3/mult_19/SUMB[7][2] ), .B(\U3/mult_19/CARRYB[7][1] ), .Q(
        \U3/mult_19/A1[7] ) );
  NOR21 U254 ( .A(\U2/n278 ), .B(n232), .Q(\U2/n738 ) );
  NOR21 U255 ( .A(\U2/n278 ), .B(Rom_Address[2]), .Q(\U2/n733 ) );
  INV3 U256 ( .A(\U2/n727 ), .Q(\U2/n266 ) );
  INV3 U257 ( .A(\U2/n726 ), .Q(\U2/n267 ) );
  INV3 U258 ( .A(\U2/n740 ), .Q(\U2/n271 ) );
  NAND22 U259 ( .A(\U2/n738 ), .B(\U2/n718 ), .Q(\U2/n740 ) );
  NOR21 U260 ( .A(\U1/n20 ), .B(n233), .Q(\U1/n24 ) );
  NOR21 U261 ( .A(\U1/n2 ), .B(n233), .Q(\U1/n17 ) );
  AOI211 U262 ( .A(\U1/n15 ), .B(\U1/n7 ), .C(\U1/n24 ), .Q(\U1/n31 ) );
  INV3 U263 ( .A(\U2/n736 ), .Q(\U2/n274 ) );
  NAND22 U264 ( .A(\U2/n733 ), .B(\U2/n717 ), .Q(\U2/n736 ) );
  INV3 U265 ( .A(\U2/n735 ), .Q(\U2/n275 ) );
  NAND22 U266 ( .A(\U2/n733 ), .B(\U2/n718 ), .Q(\U2/n735 ) );
  NAND22 U267 ( .A(\U2/n716 ), .B(\U2/n718 ), .Q(\U2/n356 ) );
  INV3 U268 ( .A(\U1/n37 ), .Q(Rom_out[7]) );
  INV3 U269 ( .A(\U3/mult_19/ab[0][5] ), .Q(\U3/mult_19/n80 ) );
  INV3 U270 ( .A(\U3/mult_19/ab[0][3] ), .Q(\U3/mult_19/n78 ) );
  INV3 U271 ( .A(\U3/mult_19/ab[1][4] ), .Q(\U3/mult_19/n72 ) );
  INV3 U272 ( .A(\U3/mult_19/ab[1][3] ), .Q(\U3/mult_19/n71 ) );
  INV3 U273 ( .A(Rom_out[0]), .Q(\U3/mult_19/n91 ) );
  OAI2111 U274 ( .A(\U1/n18 ), .B(\U1/n4 ), .C(\U1/n11 ), .D(\U1/n52 ), .Q(
        Rom_out[0]) );
  INV3 U275 ( .A(\U1/n24 ), .Q(\U1/n4 ) );
  AOI311 U276 ( .A(\U1/n16 ), .B(\U1/n7 ), .C(\U1/n15 ), .D(\U1/n53 ), .Q(
        \U1/n52 ) );
  XOR21 U277 ( .A(\U3/mult_19/SUMB[7][4] ), .B(\U3/mult_19/CARRYB[7][3] ), .Q(
        \U3/mult_19/A1[9] ) );
  XOR21 U278 ( .A(\U3/mult_19/SUMB[7][5] ), .B(\U3/mult_19/CARRYB[7][4] ), .Q(
        \U3/mult_19/A1[10] ) );
  INV3 U279 ( .A(Rom_out[2]), .Q(\U3/mult_19/n89 ) );
  NAND22 U280 ( .A(\U1/n41 ), .B(\U1/n42 ), .Q(Rom_out[2]) );
  AOI221 U281 ( .A(\U1/n44 ), .B(\U1/n2 ), .C(n233), .D(\U1/n45 ), .Q(\U1/n41 ) );
  AOI311 U282 ( .A(n232), .B(\U1/n7 ), .C(\U1/n11 ), .D(\U1/n43 ), .Q(\U1/n42 ) );
  NAND22 U283 ( .A(\U1/n9 ), .B(\U1/n7 ), .Q(\U1/n16 ) );
  NOR21 U284 ( .A(\U1/n19 ), .B(\U1/n7 ), .Q(\U1/n35 ) );
  NOR21 U285 ( .A(\U3/mult_19/n51 ), .B(\U3/mult_19/n54 ), .Q(
        \U3/mult_19/A2[9] ) );
  INV3 U286 ( .A(\U3/mult_19/CARRYB[7][2] ), .Q(\U3/mult_19/n51 ) );
  INV3 U287 ( .A(\U3/mult_19/SUMB[7][3] ), .Q(\U3/mult_19/n54 ) );
  NOR31 U288 ( .A(\U1/n3 ), .B(\U1/n28 ), .C(\U1/n35 ), .Q(\U1/n53 ) );
  INV3 U289 ( .A(\U1/n25 ), .Q(\U1/n3 ) );
  BUF2 U290 ( .A(\U2/n359 ), .Q(n236) );
  INV3 U291 ( .A(\U1/n19 ), .Q(\U1/n9 ) );
  INV3 U292 ( .A(\U1/n18 ), .Q(\U1/n5 ) );
  XOR21 U293 ( .A(\U3/mult_19/SUMB[7][6] ), .B(\U3/mult_19/CARRYB[7][5] ), .Q(
        \U3/mult_19/A1[11] ) );
  INV3 U294 ( .A(Mult_out[0]), .Q(\U4/add_27_aco/n20 ) );
  XOR21 U295 ( .A(\U3/mult_19/ab[7][7] ), .B(\U3/mult_19/CARRYB[7][6] ), .Q(
        \U3/mult_19/A1[12] ) );
  BUF2 U296 ( .A(\U2/n286 ), .Q(n250) );
  BUF2 U297 ( .A(\U2/n286 ), .Q(n249) );
  BUF2 U298 ( .A(\U2/n285 ), .Q(n245) );
  BUF2 U299 ( .A(\U2/n285 ), .Q(n248) );
  BUF2 U300 ( .A(\U2/n285 ), .Q(n246) );
  BUF2 U301 ( .A(n246), .Q(n247) );
  INV3 U302 ( .A(Rom_out[5]), .Q(\U3/mult_19/n86 ) );
  OAI2111 U303 ( .A(\U1/n19 ), .B(\U1/n20 ), .C(\U1/n21 ), .D(\U1/n22 ), .Q(
        Rom_out[5]) );
  INV3 U304 ( .A(Rom_out[6]), .Q(\U3/mult_19/n85 ) );
  NAND22 U305 ( .A(\U1/n13 ), .B(\U1/n14 ), .Q(Rom_out[6]) );
  AOI221 U306 ( .A(\U1/n18 ), .B(\U1/n2 ), .C(\U1/n6 ), .D(Rom_Address[4]), 
        .Q(\U1/n13 ) );
  AOI221 U307 ( .A(\U1/n15 ), .B(\U1/n16 ), .C(\U1/n17 ), .D(\U1/n5 ), .Q(
        \U1/n14 ) );
  XNR21 U308 ( .A(Rom_Address[4]), .B(n233), .Q(\U1/n25 ) );
  NOR21 U309 ( .A(\U2/n280 ), .B(n230), .Q(\U2/n717 ) );
  NOR21 U310 ( .A(\U2/n280 ), .B(\U1/n12 ), .Q(\U2/n718 ) );
  NOR21 U311 ( .A(\U3/mult_19/n62 ), .B(\U3/mult_19/n91 ), .Q(
        \U3/mult_19/ab[7][0] ) );
  NOR21 U312 ( .A(\U3/mult_19/n62 ), .B(\U3/mult_19/n90 ), .Q(
        \U3/mult_19/ab[7][1] ) );
  NOR21 U313 ( .A(n233), .B(n231), .Q(\U2/n724 ) );
  NOR21 U314 ( .A(\U3/mult_19/n62 ), .B(\U3/mult_19/n89 ), .Q(
        \U3/mult_19/ab[7][2] ) );
  NOR21 U315 ( .A(\U3/mult_19/n62 ), .B(\U3/mult_19/n88 ), .Q(
        \U3/mult_19/ab[7][3] ) );
  INV3 U316 ( .A(Rom_out[4]), .Q(\U3/mult_19/n87 ) );
  OAI2111 U317 ( .A(\U1/n31 ), .B(\U1/n32 ), .C(\U1/n33 ), .D(\U1/n34 ), .Q(
        Rom_out[4]) );
  NAND22 U318 ( .A(\U1/n35 ), .B(\U1/n15 ), .Q(\U1/n33 ) );
  AOI221 U319 ( .A(\U1/n28 ), .B(\U1/n17 ), .C(\U1/n25 ), .D(\U1/n32 ), .Q(
        \U1/n34 ) );
  INV3 U320 ( .A(\U2/n732 ), .Q(\U2/n277 ) );
  NAND22 U321 ( .A(\U2/n733 ), .B(\U2/n720 ), .Q(\U2/n732 ) );
  INV3 U322 ( .A(Rom_Address[4]), .Q(\U1/n2 ) );
  NOR21 U323 ( .A(\U3/mult_19/n91 ), .B(\U3/mult_19/n65 ), .Q(
        \U3/mult_19/ab[4][0] ) );
  NOR21 U324 ( .A(\U3/mult_19/n90 ), .B(\U3/mult_19/n65 ), .Q(
        \U3/mult_19/ab[4][1] ) );
  NOR21 U325 ( .A(\U3/mult_19/n89 ), .B(\U3/mult_19/n65 ), .Q(
        \U3/mult_19/ab[4][2] ) );
  NOR21 U326 ( .A(\U3/mult_19/n88 ), .B(\U3/mult_19/n65 ), .Q(
        \U3/mult_19/ab[4][3] ) );
  NOR21 U327 ( .A(\U3/mult_19/n87 ), .B(\U3/mult_19/n65 ), .Q(
        \U3/mult_19/ab[4][4] ) );
  NOR21 U328 ( .A(\U3/mult_19/n91 ), .B(\U3/mult_19/n64 ), .Q(
        \U3/mult_19/ab[5][0] ) );
  NOR21 U329 ( .A(\U3/mult_19/n90 ), .B(\U3/mult_19/n64 ), .Q(
        \U3/mult_19/ab[5][1] ) );
  NOR21 U330 ( .A(\U3/mult_19/n89 ), .B(\U3/mult_19/n64 ), .Q(
        \U3/mult_19/ab[5][2] ) );
  NOR21 U331 ( .A(\U3/mult_19/n88 ), .B(\U3/mult_19/n64 ), .Q(
        \U3/mult_19/ab[5][3] ) );
  NOR21 U332 ( .A(\U3/mult_19/n91 ), .B(\U3/mult_19/n63 ), .Q(
        \U3/mult_19/ab[6][0] ) );
  NOR21 U333 ( .A(\U3/mult_19/n90 ), .B(\U3/mult_19/n63 ), .Q(
        \U3/mult_19/ab[6][1] ) );
  NOR21 U334 ( .A(\U3/mult_19/n89 ), .B(\U3/mult_19/n63 ), .Q(
        \U3/mult_19/ab[6][2] ) );
  NOR21 U335 ( .A(\U3/mult_19/n88 ), .B(\U3/mult_19/n63 ), .Q(
        \U3/mult_19/ab[6][3] ) );
  NOR21 U336 ( .A(\U3/mult_19/n90 ), .B(\U3/mult_19/n66 ), .Q(
        \U3/mult_19/ab[3][1] ) );
  NOR21 U337 ( .A(\U3/mult_19/n89 ), .B(\U3/mult_19/n66 ), .Q(
        \U3/mult_19/ab[3][2] ) );
  NOR21 U338 ( .A(\U3/mult_19/n88 ), .B(\U3/mult_19/n66 ), .Q(
        \U3/mult_19/ab[3][3] ) );
  NOR21 U339 ( .A(\U3/mult_19/n87 ), .B(\U3/mult_19/n66 ), .Q(
        \U3/mult_19/ab[3][4] ) );
  NOR21 U340 ( .A(\U3/mult_19/n86 ), .B(\U3/mult_19/n66 ), .Q(
        \U3/mult_19/ab[3][5] ) );
  NOR21 U341 ( .A(\U3/mult_19/n90 ), .B(\U3/mult_19/n67 ), .Q(
        \U3/mult_19/ab[2][1] ) );
  XOR21 U342 ( .A(\U3/mult_19/ab[0][3] ), .B(\U3/mult_19/ab[1][2] ), .Q(
        \U3/mult_19/SUMB[1][2] ) );
  NOR21 U343 ( .A(\U3/mult_19/n89 ), .B(\U3/mult_19/n67 ), .Q(
        \U3/mult_19/ab[2][2] ) );
  NOR21 U344 ( .A(\U3/mult_19/n78 ), .B(\U3/mult_19/n70 ), .Q(
        \U3/mult_19/CARRYB[1][2] ) );
  XOR21 U345 ( .A(\U3/mult_19/ab[0][4] ), .B(\U3/mult_19/ab[1][3] ), .Q(
        \U3/mult_19/SUMB[1][3] ) );
  NOR21 U346 ( .A(\U3/mult_19/n88 ), .B(\U3/mult_19/n67 ), .Q(
        \U3/mult_19/ab[2][3] ) );
  NOR21 U347 ( .A(\U3/mult_19/n79 ), .B(\U3/mult_19/n71 ), .Q(
        \U3/mult_19/CARRYB[1][3] ) );
  XOR21 U348 ( .A(\U3/mult_19/ab[0][5] ), .B(\U3/mult_19/ab[1][4] ), .Q(
        \U3/mult_19/SUMB[1][4] ) );
  NOR21 U349 ( .A(\U3/mult_19/n87 ), .B(\U3/mult_19/n67 ), .Q(
        \U3/mult_19/ab[2][4] ) );
  NOR21 U350 ( .A(\U3/mult_19/n80 ), .B(\U3/mult_19/n72 ), .Q(
        \U3/mult_19/CARRYB[1][4] ) );
  XOR21 U351 ( .A(\U3/mult_19/ab[0][6] ), .B(\U3/mult_19/ab[1][5] ), .Q(
        \U3/mult_19/SUMB[1][5] ) );
  NOR21 U352 ( .A(\U3/mult_19/n86 ), .B(\U3/mult_19/n67 ), .Q(
        \U3/mult_19/ab[2][5] ) );
  XOR21 U353 ( .A(\U3/mult_19/ab[0][7] ), .B(\U3/mult_19/ab[1][6] ), .Q(
        \U3/mult_19/SUMB[1][6] ) );
  NOR21 U354 ( .A(\U3/mult_19/n87 ), .B(\U3/mult_19/n75 ), .Q(
        \U3/mult_19/ab[1][4] ) );
  NOR21 U355 ( .A(\U3/mult_19/n86 ), .B(\U3/mult_19/n75 ), .Q(
        \U3/mult_19/ab[1][5] ) );
  NOR21 U356 ( .A(\U3/mult_19/n85 ), .B(\U3/mult_19/n75 ), .Q(
        \U3/mult_19/ab[1][6] ) );
  NOR21 U357 ( .A(\U3/mult_19/n86 ), .B(\U3/mult_19/n83 ), .Q(
        \U3/mult_19/ab[0][5] ) );
  NOR21 U358 ( .A(\U3/mult_19/n85 ), .B(\U3/mult_19/n83 ), .Q(
        \U3/mult_19/ab[0][6] ) );
  NOR21 U359 ( .A(\U3/mult_19/n84 ), .B(\U3/mult_19/n83 ), .Q(
        \U3/mult_19/ab[0][7] ) );
  INV3 U360 ( .A(\U2/n739 ), .Q(\U2/n272 ) );
  NAND22 U361 ( .A(\U2/n738 ), .B(\U2/n719 ), .Q(\U2/n739 ) );
  NOR21 U362 ( .A(\U3/mult_19/n84 ), .B(\U3/mult_19/n67 ), .Q(
        \U3/mult_19/ab[2][7] ) );
  NOR21 U363 ( .A(\U3/mult_19/n85 ), .B(\U3/mult_19/n66 ), .Q(
        \U3/mult_19/ab[3][6] ) );
  NOR21 U364 ( .A(\U3/mult_19/n86 ), .B(\U3/mult_19/n65 ), .Q(
        \U3/mult_19/ab[4][5] ) );
  NOR21 U365 ( .A(\U3/mult_19/n84 ), .B(\U3/mult_19/n66 ), .Q(
        \U3/mult_19/ab[3][7] ) );
  NOR21 U366 ( .A(\U3/mult_19/n85 ), .B(\U3/mult_19/n65 ), .Q(
        \U3/mult_19/ab[4][6] ) );
  NOR21 U367 ( .A(\U3/mult_19/n87 ), .B(\U3/mult_19/n64 ), .Q(
        \U3/mult_19/ab[5][4] ) );
  NOR21 U368 ( .A(\U3/mult_19/n86 ), .B(\U3/mult_19/n64 ), .Q(
        \U3/mult_19/ab[5][5] ) );
  NOR21 U369 ( .A(\U3/mult_19/n87 ), .B(\U3/mult_19/n63 ), .Q(
        \U3/mult_19/ab[6][4] ) );
  INV3 U370 ( .A(n232), .Q(n233) );
  NOR21 U371 ( .A(\U3/mult_19/n85 ), .B(\U3/mult_19/n67 ), .Q(
        \U3/mult_19/ab[2][6] ) );
  INV3 U372 ( .A(Rom_out[3]), .Q(\U3/mult_19/n88 ) );
  AOI2111 U373 ( .A(\U1/n9 ), .B(\U1/n20 ), .C(\U1/n38 ), .D(\U1/n39 ), .Q(
        \U1/n36 ) );
  XNR21 U374 ( .A(\U2/n280 ), .B(n233), .Q(\U1/n38 ) );
  NOR21 U375 ( .A(\U3/mult_19/n62 ), .B(\U3/mult_19/n87 ), .Q(
        \U3/mult_19/ab[7][4] ) );
  NOR21 U376 ( .A(\U3/mult_19/n62 ), .B(\U3/mult_19/n86 ), .Q(
        \U3/mult_19/ab[7][5] ) );
  NOR21 U377 ( .A(n232), .B(Rom_Address[4]), .Q(\U1/n15 ) );
  OAI2111 U378 ( .A(\U1/n7 ), .B(\U1/n32 ), .C(\U1/n20 ), .D(\U1/n46 ), .Q(
        \U1/n45 ) );
  NAND22 U379 ( .A(Rom_Address[4]), .B(\U1/n12 ), .Q(\U1/n46 ) );
  NOR21 U380 ( .A(\U1/n40 ), .B(\U1/n7 ), .Q(\U1/n18 ) );
  NAND22 U381 ( .A(\U1/n12 ), .B(\U2/n280 ), .Q(\U1/n19 ) );
  NOR21 U382 ( .A(\U3/mult_19/n91 ), .B(\U3/mult_19/n66 ), .Q(
        \U3/mult_19/ab[3][0] ) );
  NOR21 U383 ( .A(\U3/mult_19/n91 ), .B(\U3/mult_19/n67 ), .Q(
        \U3/mult_19/ab[2][0] ) );
  XOR21 U384 ( .A(\U3/mult_19/ab[0][2] ), .B(\U3/mult_19/ab[1][1] ), .Q(
        \U3/mult_19/SUMB[1][1] ) );
  AOI211 U385 ( .A(\U1/n29 ), .B(\U1/n30 ), .C(\U1/n7 ), .Q(\U1/n27 ) );
  INV3 U386 ( .A(Rom_out[1]), .Q(\U3/mult_19/n90 ) );
  AOI221 U387 ( .A(n233), .B(\U1/n50 ), .C(\U1/n6 ), .D(\U1/n17 ), .Q(\U1/n49 ) );
  NOR21 U388 ( .A(\U3/mult_19/n84 ), .B(\U3/mult_19/n65 ), .Q(
        \U3/mult_19/ab[4][7] ) );
  NOR21 U389 ( .A(\U3/mult_19/n85 ), .B(\U3/mult_19/n64 ), .Q(
        \U3/mult_19/ab[5][6] ) );
  NOR21 U390 ( .A(\U3/mult_19/n86 ), .B(\U3/mult_19/n63 ), .Q(
        \U3/mult_19/ab[6][5] ) );
  NOR21 U391 ( .A(\U3/mult_19/n84 ), .B(\U3/mult_19/n64 ), .Q(
        \U3/mult_19/ab[5][7] ) );
  NOR21 U392 ( .A(\U3/mult_19/n85 ), .B(\U3/mult_19/n63 ), .Q(
        \U3/mult_19/ab[6][6] ) );
  INV3 U393 ( .A(\U1/n32 ), .Q(\U1/n11 ) );
  NOR21 U394 ( .A(\U1/n40 ), .B(\U1/n20 ), .Q(\U1/n39 ) );
  NOR21 U395 ( .A(\U3/mult_19/n84 ), .B(\U3/mult_19/n63 ), .Q(
        \U3/mult_19/ab[6][7] ) );
  NOR21 U396 ( .A(\U3/mult_19/n62 ), .B(\U3/mult_19/n85 ), .Q(
        \U3/mult_19/ab[7][6] ) );
  NOR21 U397 ( .A(\U3/mult_19/n62 ), .B(\U3/mult_19/n84 ), .Q(
        \U3/mult_19/ab[7][7] ) );
  NOR21 U398 ( .A(RESET), .B(\U4/n42 ), .Q(\U4/N28 ) );
  INV3 U399 ( .A(\U4/N7 ), .Q(\U4/n42 ) );
  NOR21 U400 ( .A(RESET), .B(\U2/n285 ), .Q(\U2/n286 ) );
  INV3 U401 ( .A(\U6/n28 ), .Q(\U6/n7 ) );
  NOR22 U402 ( .A(\U5/n11 ), .B(RESET), .Q(\U5/n3 ) );
  INV3 U403 ( .A(\U5/n11 ), .Q(\U5/n1 ) );
  INV3 U404 ( .A(\U8/n5 ), .Q(\U8/n1 ) );
  NOR21 U405 ( .A(n230), .B(n229), .Q(\U2/n719 ) );
  NOR21 U406 ( .A(\U1/n12 ), .B(n229), .Q(\U2/n720 ) );
  INV3 U407 ( .A(\U6/n29 ), .Q(Rom_Address[4]) );
  NOR40 U408 ( .A(\U2/n712 ), .B(\U2/n713 ), .C(\U2/n714 ), .D(\U2/n715 ), .Q(
        \U2/n700 ) );
  NOR40 U409 ( .A(\U2/n702 ), .B(\U2/n703 ), .C(\U2/n704 ), .D(\U2/n705 ), .Q(
        \U2/n701 ) );
  INV3 U410 ( .A(Delay_Line_out[2]), .Q(\U3/mult_19/n67 ) );
  NOR40 U411 ( .A(\U2/n668 ), .B(\U2/n669 ), .C(\U2/n670 ), .D(\U2/n671 ), .Q(
        \U2/n656 ) );
  NOR40 U412 ( .A(\U2/n658 ), .B(\U2/n659 ), .C(\U2/n660 ), .D(\U2/n661 ), .Q(
        \U2/n657 ) );
  NOR40 U413 ( .A(\U2/n690 ), .B(\U2/n691 ), .C(\U2/n692 ), .D(\U2/n693 ), .Q(
        \U2/n678 ) );
  NOR40 U414 ( .A(\U2/n680 ), .B(\U2/n681 ), .C(\U2/n682 ), .D(\U2/n683 ), .Q(
        \U2/n679 ) );
  INV3 U415 ( .A(Delay_Line_out[3]), .Q(\U3/mult_19/n66 ) );
  NOR40 U416 ( .A(\U2/n646 ), .B(\U2/n647 ), .C(\U2/n648 ), .D(\U2/n649 ), .Q(
        \U2/n634 ) );
  NOR40 U417 ( .A(\U2/n636 ), .B(\U2/n637 ), .C(\U2/n638 ), .D(\U2/n639 ), .Q(
        \U2/n635 ) );
  NOR21 U418 ( .A(RESET), .B(n224), .Q(\U4/N46 ) );
  INV3 U419 ( .A(\U6/n44 ), .Q(\U6/n11 ) );
  INV3 U420 ( .A(Rom_Address[2]), .Q(n232) );
  NOR21 U421 ( .A(n19), .B(\U6/n44 ), .Q(Rom_Address[2]) );
  BUF2 U422 ( .A(Rom_Address[3]), .Q(n231) );
  NOR21 U423 ( .A(n31), .B(\U6/n44 ), .Q(Rom_Address[3]) );
  NOR21 U424 ( .A(\U4/add_27_aco/n14 ), .B(\U4/mult_add_27_aco/PROD_not[18] ), 
        .Q(\U4/add_27_aco/carry [19]) );
  INV3 U425 ( .A(\U4/add_27_aco/carry [18]), .Q(\U4/add_27_aco/n14 ) );
  NOR21 U426 ( .A(\U4/add_27_aco/n18 ), .B(\U4/mult_add_27_aco/PROD_not[16] ), 
        .Q(\U4/add_27_aco/carry [17]) );
  NOR40 U427 ( .A(\U2/n624 ), .B(\U2/n625 ), .C(\U2/n626 ), .D(\U2/n627 ), .Q(
        \U2/n612 ) );
  NOR40 U428 ( .A(\U2/n614 ), .B(\U2/n615 ), .C(\U2/n616 ), .D(\U2/n617 ), .Q(
        \U2/n613 ) );
  INV3 U429 ( .A(\U4/mult_add_27_aco/PROD_not[1] ), .Q(\U4/N49 ) );
  NOR21 U430 ( .A(\U4/add_27_aco/n20 ), .B(\U4/mult_add_27_aco/PROD_not[0] ), 
        .Q(\U4/add_27_aco/carry [1]) );
  XOR21 U431 ( .A(\U3/mult_19/ab[0][1] ), .B(\U3/mult_19/ab[1][0] ), .Q(
        Mult_out[1]) );
  NOR21 U432 ( .A(RESET), .B(\U4/n29 ), .Q(\U4/N41 ) );
  INV3 U433 ( .A(\U4/N20 ), .Q(\U4/n29 ) );
  NOR21 U434 ( .A(RESET), .B(\U4/n28 ), .Q(\U4/N42 ) );
  INV3 U435 ( .A(\U4/N21 ), .Q(\U4/n28 ) );
  NOR40 U436 ( .A(\U2/n602 ), .B(\U2/n603 ), .C(\U2/n604 ), .D(\U2/n605 ), .Q(
        \U2/n522 ) );
  NOR40 U437 ( .A(\U2/n592 ), .B(\U2/n593 ), .C(\U2/n594 ), .D(\U2/n595 ), .Q(
        \U2/n523 ) );
  INV3 U438 ( .A(Delay_Line_out[6]), .Q(\U3/mult_19/n63 ) );
  NOR40 U439 ( .A(\U2/n388 ), .B(\U2/n389 ), .C(\U2/n390 ), .D(\U2/n391 ), .Q(
        \U2/n376 ) );
  NOR40 U440 ( .A(\U2/n378 ), .B(\U2/n379 ), .C(\U2/n380 ), .D(\U2/n381 ), .Q(
        \U2/n377 ) );
  NOR21 U441 ( .A(RESET), .B(\U4/n30 ), .Q(\U4/N40 ) );
  INV3 U442 ( .A(\U4/N19 ), .Q(\U4/n30 ) );
  NOR21 U443 ( .A(RESET), .B(\U4/n31 ), .Q(\U4/N39 ) );
  INV3 U444 ( .A(\U4/N18 ), .Q(\U4/n31 ) );
  NOR21 U445 ( .A(RESET), .B(\U4/n32 ), .Q(\U4/N38 ) );
  INV3 U446 ( .A(\U4/N17 ), .Q(\U4/n32 ) );
  NOR40 U447 ( .A(\U2/n366 ), .B(\U2/n367 ), .C(\U2/n368 ), .D(\U2/n369 ), .Q(
        \U2/n350 ) );
  NOR40 U448 ( .A(\U2/n352 ), .B(\U2/n353 ), .C(\U2/n354 ), .D(\U2/n355 ), .Q(
        \U2/n351 ) );
  NOR21 U449 ( .A(RESET), .B(\U4/n33 ), .Q(\U4/N37 ) );
  INV3 U450 ( .A(\U4/N16 ), .Q(\U4/n33 ) );
  BUF2 U451 ( .A(\U6/n24 ), .Q(n234) );
  NOR21 U452 ( .A(RESET), .B(\U4/n35 ), .Q(\U4/N35 ) );
  INV3 U453 ( .A(\U4/N14 ), .Q(\U4/n35 ) );
  NOR21 U454 ( .A(RESET), .B(\U4/n34 ), .Q(\U4/N36 ) );
  INV3 U455 ( .A(\U4/N15 ), .Q(\U4/n34 ) );
  NOR21 U456 ( .A(RESET), .B(\U4/n36 ), .Q(\U4/N34 ) );
  INV3 U457 ( .A(\U4/N13 ), .Q(\U4/n36 ) );
  NOR21 U458 ( .A(RESET), .B(\U4/n37 ), .Q(\U4/N33 ) );
  INV3 U459 ( .A(\U4/N12 ), .Q(\U4/n37 ) );
  NOR21 U460 ( .A(RESET), .B(\U4/n39 ), .Q(\U4/N31 ) );
  INV3 U461 ( .A(\U4/N10 ), .Q(\U4/n39 ) );
  NOR21 U462 ( .A(RESET), .B(\U4/n38 ), .Q(\U4/N32 ) );
  INV3 U463 ( .A(\U4/N11 ), .Q(\U4/n38 ) );
  NOR21 U464 ( .A(RESET), .B(\U4/n40 ), .Q(\U4/N30 ) );
  INV3 U465 ( .A(\U4/N9 ), .Q(\U4/n40 ) );
  NOR21 U466 ( .A(RESET), .B(\U4/n41 ), .Q(\U4/N29 ) );
  INV3 U467 ( .A(\U4/N8 ), .Q(\U4/n41 ) );
  INV3 U468 ( .A(ack_F2ADC), .Q(\U6/n16 ) );
  NOR21 U469 ( .A(RESET), .B(Delay_Line_sample_shift), .Q(\U2/n285 ) );
  OAI2111 U470 ( .A(\U6/n27 ), .B(\U1/n7 ), .C(\U6/n32 ), .D(\U6/n34 ), .Q(
        \U6/n40 ) );
  NAND31 U471 ( .A(\U6/n11 ), .B(n31), .C(\U6/n27 ), .Q(\U6/n32 ) );
  NAND31 U472 ( .A(\U6/n16 ), .B(\U6/n28 ), .C(\U6/n46 ), .Q(\U6/n37 ) );
  AOI211 U473 ( .A(\U6/n11 ), .B(n121), .C(\U6/n31 ), .Q(\U6/n46 ) );
  NOR21 U474 ( .A(Buff_OE), .B(\U6/n8 ), .Q(\U6/n28 ) );
  INV3 U475 ( .A(\U6/n34 ), .Q(\U6/n8 ) );
  NOR22 U476 ( .A(\U9/n11 ), .B(RESET), .Q(\U9/n3 ) );
  INV3 U477 ( .A(\U9/n11 ), .Q(\U9/n1 ) );
  NOR21 U478 ( .A(Buff_OE), .B(RESET), .Q(\U5/n11 ) );
  INV3 U479 ( .A(\U6/n27 ), .Q(\U6/n13 ) );
  NAND22 U480 ( .A(req_F2DAC), .B(n263), .Q(\U8/n5 ) );
  INV3 U481 ( .A(\U6/n23 ), .Q(req_F2DAC) );
  INV3 U482 ( .A(\U7/n12 ), .Q(req_ADC2F) );
  NOR21 U483 ( .A(req_ADC2F), .B(\U7/n1 ), .Q(\U7/n14 ) );
  INV3 U484 ( .A(ADC_Rdb), .Q(\U7/n1 ) );
  INV3 U485 ( .A(\U4/mult_add_27_aco/PROD_not[15] ), .Q(\U4/N63 ) );
  NAND22 U486 ( .A(Accu_out[15]), .B(\U6/n24 ), .Q(
        \U4/mult_add_27_aco/PROD_not[15] ) );
  NAND41 U487 ( .A(\U2/n708 ), .B(\U2/n709 ), .C(\U2/n710 ), .D(\U2/n711 ), 
        .Q(\U2/n702 ) );
  AOI221 U488 ( .A(\U2/n274 ), .B(\U2/x[26][0] ), .C(\U2/n275 ), .D(
        \U2/x[27][0] ), .Q(\U2/n710 ) );
  AOI221 U489 ( .A(\U2/n276 ), .B(\U2/x[24][0] ), .C(\U2/n277 ), .D(
        \U2/x[25][0] ), .Q(\U2/n711 ) );
  AOI221 U490 ( .A(\U2/n270 ), .B(\U2/x[30][0] ), .C(\U2/n271 ), .D(
        \U2/x[31][0] ), .Q(\U2/n708 ) );
  NAND41 U491 ( .A(\U2/n728 ), .B(\U2/n729 ), .C(\U2/n730 ), .D(\U2/n731 ), 
        .Q(\U2/n712 ) );
  NAND41 U492 ( .A(\U2/n664 ), .B(\U2/n665 ), .C(\U2/n666 ), .D(\U2/n667 ), 
        .Q(\U2/n658 ) );
  NAND41 U493 ( .A(\U2/n674 ), .B(\U2/n675 ), .C(\U2/n676 ), .D(\U2/n677 ), 
        .Q(\U2/n668 ) );
  NAND41 U494 ( .A(\U2/n686 ), .B(\U2/n687 ), .C(\U2/n688 ), .D(\U2/n689 ), 
        .Q(\U2/n680 ) );
  AOI221 U495 ( .A(\U2/n274 ), .B(\U2/x[26][1] ), .C(\U2/n275 ), .D(
        \U2/x[27][1] ), .Q(\U2/n688 ) );
  AOI221 U496 ( .A(\U2/n276 ), .B(\U2/x[24][1] ), .C(\U2/n277 ), .D(
        \U2/x[25][1] ), .Q(\U2/n689 ) );
  AOI221 U497 ( .A(\U2/n270 ), .B(\U2/x[30][1] ), .C(\U2/n271 ), .D(
        \U2/x[31][1] ), .Q(\U2/n686 ) );
  NAND41 U498 ( .A(\U2/n696 ), .B(\U2/n697 ), .C(\U2/n698 ), .D(\U2/n699 ), 
        .Q(\U2/n690 ) );
  NAND41 U499 ( .A(\U2/n642 ), .B(\U2/n643 ), .C(\U2/n644 ), .D(\U2/n645 ), 
        .Q(\U2/n636 ) );
  NAND22 U500 ( .A(\U6/n48 ), .B(\U6/n11 ), .Q(\U6/n29 ) );
  AOI221 U501 ( .A(\U2/n272 ), .B(\U2/x[28][0] ), .C(\U2/n273 ), .D(
        \U2/x[29][0] ), .Q(\U2/n709 ) );
  AOI221 U502 ( .A(\U2/n272 ), .B(\U2/x[28][1] ), .C(\U2/n273 ), .D(
        \U2/x[29][1] ), .Q(\U2/n687 ) );
  INV3 U503 ( .A(\U4/mult_add_27_aco/PROD_not[14] ), .Q(\U4/N62 ) );
  NAND22 U504 ( .A(Accu_out[14]), .B(n234), .Q(
        \U4/mult_add_27_aco/PROD_not[14] ) );
  INV3 U505 ( .A(\U4/mult_add_27_aco/PROD_not[10] ), .Q(\U4/N58 ) );
  NAND22 U506 ( .A(\U4/Accu_out[10] ), .B(n234), .Q(
        \U4/mult_add_27_aco/PROD_not[10] ) );
  INV3 U507 ( .A(\U4/mult_add_27_aco/PROD_not[8] ), .Q(\U4/N56 ) );
  NAND22 U508 ( .A(\U4/Accu_out[8] ), .B(\U6/n24 ), .Q(
        \U4/mult_add_27_aco/PROD_not[8] ) );
  INV3 U509 ( .A(\U4/mult_add_27_aco/PROD_not[12] ), .Q(\U4/N60 ) );
  NAND22 U510 ( .A(Accu_out[12]), .B(n234), .Q(
        \U4/mult_add_27_aco/PROD_not[12] ) );
  INV3 U511 ( .A(\U4/mult_add_27_aco/PROD_not[9] ), .Q(\U4/N57 ) );
  NAND22 U512 ( .A(n234), .B(\U4/Accu_out[9] ), .Q(
        \U4/mult_add_27_aco/PROD_not[9] ) );
  INV3 U513 ( .A(\U4/mult_add_27_aco/PROD_not[11] ), .Q(\U4/N59 ) );
  XNR21 U514 ( .A(\U3/mult_19/FS_1/n9 ), .B(\U3/mult_19/FS_1/n10 ), .Q(
        Mult_out[11]) );
  NAND22 U515 ( .A(\U4/Accu_out[11] ), .B(\U6/n24 ), .Q(
        \U4/mult_add_27_aco/PROD_not[11] ) );
  INV3 U516 ( .A(\U4/mult_add_27_aco/PROD_not[6] ), .Q(\U4/N54 ) );
  NAND22 U517 ( .A(\U4/Accu_out[6] ), .B(n234), .Q(
        \U4/mult_add_27_aco/PROD_not[6] ) );
  INV3 U518 ( .A(\U4/mult_add_27_aco/PROD_not[7] ), .Q(\U4/N55 ) );
  NAND22 U519 ( .A(\U4/Accu_out[7] ), .B(n234), .Q(
        \U4/mult_add_27_aco/PROD_not[7] ) );
  NAND22 U520 ( .A(\U2/n706 ), .B(\U2/n707 ), .Q(\U2/n703 ) );
  AOI221 U521 ( .A(\U2/n266 ), .B(\U2/x[18][0] ), .C(\U2/n267 ), .D(
        \U2/x[19][0] ), .Q(\U2/n706 ) );
  AOI221 U522 ( .A(\U2/n268 ), .B(\U2/x[16][0] ), .C(\U2/n269 ), .D(
        \U2/x[17][0] ), .Q(\U2/n707 ) );
  NAND22 U523 ( .A(\U2/n721 ), .B(\U2/n722 ), .Q(\U2/n713 ) );
  AOI221 U524 ( .A(\U2/n266 ), .B(\U2/x[2][0] ), .C(\U2/n267 ), .D(
        \U2/x[3][0] ), .Q(\U2/n721 ) );
  NAND22 U525 ( .A(\U2/n662 ), .B(\U2/n663 ), .Q(\U2/n659 ) );
  NAND22 U526 ( .A(\U2/n672 ), .B(\U2/n673 ), .Q(\U2/n669 ) );
  NAND22 U527 ( .A(\U2/n684 ), .B(\U2/n685 ), .Q(\U2/n681 ) );
  AOI221 U528 ( .A(\U2/n266 ), .B(\U2/x[18][1] ), .C(\U2/n267 ), .D(
        \U2/x[19][1] ), .Q(\U2/n684 ) );
  AOI221 U529 ( .A(\U2/n268 ), .B(\U2/x[16][1] ), .C(\U2/n269 ), .D(
        \U2/x[17][1] ), .Q(\U2/n685 ) );
  NAND22 U530 ( .A(\U2/n694 ), .B(\U2/n695 ), .Q(\U2/n691 ) );
  AOI221 U531 ( .A(\U2/n266 ), .B(\U2/x[2][1] ), .C(\U2/n267 ), .D(
        \U2/x[3][1] ), .Q(\U2/n694 ) );
  NAND41 U532 ( .A(\U2/n652 ), .B(\U2/n653 ), .C(\U2/n654 ), .D(\U2/n655 ), 
        .Q(\U2/n646 ) );
  NAND41 U533 ( .A(\U2/n620 ), .B(\U2/n621 ), .C(\U2/n622 ), .D(\U2/n623 ), 
        .Q(\U2/n614 ) );
  NAND41 U534 ( .A(\U2/n630 ), .B(\U2/n631 ), .C(\U2/n632 ), .D(\U2/n633 ), 
        .Q(\U2/n624 ) );
  INV3 U535 ( .A(\U4/mult_add_27_aco/PROD_not[2] ), .Q(\U4/N50 ) );
  NAND22 U536 ( .A(\U4/Accu_out[2] ), .B(n234), .Q(
        \U4/mult_add_27_aco/PROD_not[2] ) );
  INV3 U537 ( .A(\U4/mult_add_27_aco/PROD_not[3] ), .Q(\U4/N51 ) );
  NAND22 U538 ( .A(\U4/Accu_out[3] ), .B(n234), .Q(
        \U4/mult_add_27_aco/PROD_not[3] ) );
  INV3 U539 ( .A(\U4/mult_add_27_aco/PROD_not[4] ), .Q(\U4/N52 ) );
  NAND22 U540 ( .A(\U4/Accu_out[4] ), .B(n234), .Q(
        \U4/mult_add_27_aco/PROD_not[4] ) );
  INV3 U541 ( .A(\U4/mult_add_27_aco/PROD_not[5] ), .Q(\U4/N53 ) );
  NAND22 U542 ( .A(\U4/Accu_out[5] ), .B(n234), .Q(
        \U4/mult_add_27_aco/PROD_not[5] ) );
  NAND22 U543 ( .A(\U2/n640 ), .B(\U2/n641 ), .Q(\U2/n637 ) );
  NAND22 U544 ( .A(\U2/n650 ), .B(\U2/n651 ), .Q(\U2/n647 ) );
  NAND22 U545 ( .A(\U2/n618 ), .B(\U2/n619 ), .Q(\U2/n615 ) );
  NAND22 U546 ( .A(\U2/n628 ), .B(\U2/n629 ), .Q(\U2/n625 ) );
  NAND41 U547 ( .A(\U2/n598 ), .B(\U2/n599 ), .C(\U2/n600 ), .D(\U2/n601 ), 
        .Q(\U2/n592 ) );
  NAND41 U548 ( .A(\U2/n608 ), .B(\U2/n609 ), .C(\U2/n610 ), .D(\U2/n611 ), 
        .Q(\U2/n602 ) );
  NAND41 U549 ( .A(\U2/n384 ), .B(\U2/n385 ), .C(\U2/n386 ), .D(\U2/n387 ), 
        .Q(\U2/n378 ) );
  NAND41 U550 ( .A(\U2/n518 ), .B(\U2/n519 ), .C(\U2/n520 ), .D(\U2/n521 ), 
        .Q(\U2/n388 ) );
  NAND22 U551 ( .A(\U2/n596 ), .B(\U2/n597 ), .Q(\U2/n593 ) );
  NAND22 U552 ( .A(\U2/n606 ), .B(\U2/n607 ), .Q(\U2/n603 ) );
  NAND22 U553 ( .A(\U2/n382 ), .B(\U2/n383 ), .Q(\U2/n379 ) );
  NAND22 U554 ( .A(\U2/n516 ), .B(\U2/n517 ), .Q(\U2/n389 ) );
  NAND41 U555 ( .A(\U2/n362 ), .B(\U2/n363 ), .C(\U2/n364 ), .D(\U2/n365 ), 
        .Q(\U2/n352 ) );
  NAND41 U556 ( .A(\U2/n372 ), .B(\U2/n373 ), .C(\U2/n374 ), .D(\U2/n375 ), 
        .Q(\U2/n366 ) );
  NAND22 U557 ( .A(\U2/n360 ), .B(\U2/n361 ), .Q(\U2/n353 ) );
  NAND22 U558 ( .A(\U2/n370 ), .B(\U2/n371 ), .Q(\U2/n367 ) );
  NOR21 U559 ( .A(\U6/n14 ), .B(\U6/n50 ), .Q(ack_F2ADC) );
  NAND22 U560 ( .A(\U4/Accu_out[1] ), .B(n234), .Q(
        \U4/mult_add_27_aco/PROD_not[1] ) );
  NAND22 U561 ( .A(\U4/Accu_out[0] ), .B(\U6/n24 ), .Q(
        \U4/mult_add_27_aco/PROD_not[0] ) );
  NAND22 U562 ( .A(\U6/n2 ), .B(ack_F2ADC), .Q(\U6/n24 ) );
  NAND31 U563 ( .A(\U6/n47 ), .B(\U6/n27 ), .C(Rom_Address[4]), .Q(\U6/n34 )
         );
  OAI2111 U564 ( .A(\U1/n12 ), .B(n223), .C(\U6/n34 ), .D(\U6/n43 ), .Q(
        \U6/n38 ) );
  INV3 U565 ( .A(\U2/n287 ), .Q(\U2/n3 ) );
  AOI221 U566 ( .A(n248), .B(\U2/x[1][6] ), .C(n250), .D(\U2/x[0][6] ), .Q(
        \U2/n287 ) );
  INV3 U567 ( .A(\U2/n288 ), .Q(\U2/n5 ) );
  AOI221 U568 ( .A(n248), .B(\U2/x[1][5] ), .C(n261), .D(\U2/x[0][5] ), .Q(
        \U2/n288 ) );
  NAND31 U569 ( .A(\U6/n35 ), .B(\U6/n34 ), .C(\U6/n36 ), .Q(\U6/n39 ) );
  INV3 U570 ( .A(\U4/mult_add_27_aco/PROD_not[16] ), .Q(\U4/N64 ) );
  NAND22 U571 ( .A(Accu_out[16]), .B(n234), .Q(
        \U4/mult_add_27_aco/PROD_not[16] ) );
  INV3 U572 ( .A(\U4/mult_add_27_aco/PROD_not[17] ), .Q(\U4/N65 ) );
  NAND22 U573 ( .A(Accu_out[17]), .B(\U6/n24 ), .Q(
        \U4/mult_add_27_aco/PROD_not[17] ) );
  INV3 U574 ( .A(\U4/mult_add_27_aco/PROD_not[18] ), .Q(\U4/N66 ) );
  NAND22 U575 ( .A(Accu_out[18]), .B(n234), .Q(
        \U4/mult_add_27_aco/PROD_not[18] ) );
  INV3 U576 ( .A(\U2/n349 ), .Q(\U2/n2 ) );
  AOI221 U577 ( .A(\U2/x[0][7] ), .B(\U2/n285 ), .C(n261), .D(Filter_In_mem[7]), .Q(\U2/n349 ) );
  INV3 U578 ( .A(\U2/n302 ), .Q(\U2/n25 ) );
  AOI221 U579 ( .A(n246), .B(\U2/x[3][7] ), .C(\U2/n286 ), .D(\U2/x[2][7] ), 
        .Q(\U2/n302 ) );
  INV3 U580 ( .A(\U2/n303 ), .Q(\U2/n26 ) );
  AOI221 U581 ( .A(n248), .B(\U2/x[3][6] ), .C(n262), .D(\U2/x[2][6] ), .Q(
        \U2/n303 ) );
  INV3 U582 ( .A(\U2/n304 ), .Q(\U2/n27 ) );
  AOI221 U583 ( .A(n248), .B(\U2/x[3][5] ), .C(n261), .D(\U2/x[2][5] ), .Q(
        \U2/n304 ) );
  INV3 U584 ( .A(\U2/n305 ), .Q(\U2/n28 ) );
  AOI221 U585 ( .A(n247), .B(\U2/x[3][4] ), .C(\U2/n286 ), .D(\U2/x[2][4] ), 
        .Q(\U2/n305 ) );
  INV3 U586 ( .A(\U2/n306 ), .Q(\U2/n29 ) );
  AOI221 U587 ( .A(n246), .B(\U2/x[3][3] ), .C(\U2/n286 ), .D(\U2/x[2][3] ), 
        .Q(\U2/n306 ) );
  INV3 U588 ( .A(\U2/n307 ), .Q(\U2/n30 ) );
  AOI221 U589 ( .A(n245), .B(\U2/x[3][2] ), .C(n261), .D(\U2/x[2][2] ), .Q(
        \U2/n307 ) );
  INV3 U590 ( .A(\U2/n308 ), .Q(\U2/n31 ) );
  AOI221 U591 ( .A(n246), .B(\U2/x[3][1] ), .C(n250), .D(\U2/x[2][1] ), .Q(
        \U2/n308 ) );
  INV3 U592 ( .A(\U2/n309 ), .Q(\U2/n32 ) );
  AOI221 U593 ( .A(n246), .B(\U2/x[3][0] ), .C(n262), .D(\U2/x[2][0] ), .Q(
        \U2/n309 ) );
  INV3 U594 ( .A(\U2/n348 ), .Q(\U2/n4 ) );
  AOI221 U595 ( .A(n246), .B(\U2/x[0][6] ), .C(n262), .D(Filter_In_mem[6]), 
        .Q(\U2/n348 ) );
  INV3 U596 ( .A(\U2/n347 ), .Q(\U2/n6 ) );
  AOI221 U597 ( .A(n248), .B(\U2/x[0][5] ), .C(n249), .D(Filter_In_mem[5]), 
        .Q(\U2/n347 ) );
  INV3 U598 ( .A(\U2/n346 ), .Q(\U2/n8 ) );
  AOI221 U599 ( .A(n246), .B(\U2/x[0][4] ), .C(n262), .D(Filter_In_mem[4]), 
        .Q(\U2/n346 ) );
  INV3 U600 ( .A(\U2/n345 ), .Q(\U2/n10 ) );
  AOI221 U601 ( .A(n247), .B(\U2/x[0][3] ), .C(n249), .D(Filter_In_mem[3]), 
        .Q(\U2/n345 ) );
  INV3 U602 ( .A(\U2/n344 ), .Q(\U2/n12 ) );
  AOI221 U603 ( .A(n247), .B(\U2/x[0][2] ), .C(n261), .D(Filter_In_mem[2]), 
        .Q(\U2/n344 ) );
  INV3 U604 ( .A(\U2/n343 ), .Q(\U2/n14 ) );
  AOI221 U605 ( .A(n246), .B(\U2/x[0][1] ), .C(n261), .D(Filter_In_mem[1]), 
        .Q(\U2/n343 ) );
  INV3 U606 ( .A(\U2/n342 ), .Q(\U2/n16 ) );
  AOI221 U607 ( .A(n245), .B(\U2/x[0][0] ), .C(n261), .D(Filter_In_mem[0]), 
        .Q(\U2/n342 ) );
  INV3 U608 ( .A(\U2/n284 ), .Q(\U2/n1 ) );
  AOI221 U609 ( .A(n247), .B(\U2/x[1][7] ), .C(n262), .D(\U2/x[0][7] ), .Q(
        \U2/n284 ) );
  INV3 U610 ( .A(\U2/n289 ), .Q(\U2/n7 ) );
  AOI221 U611 ( .A(n247), .B(\U2/x[1][4] ), .C(\U2/n286 ), .D(\U2/x[0][4] ), 
        .Q(\U2/n289 ) );
  INV3 U612 ( .A(\U2/n290 ), .Q(\U2/n9 ) );
  AOI221 U613 ( .A(n245), .B(\U2/x[1][3] ), .C(n250), .D(\U2/x[0][3] ), .Q(
        \U2/n290 ) );
  INV3 U614 ( .A(\U2/n291 ), .Q(\U2/n11 ) );
  AOI221 U615 ( .A(n246), .B(\U2/x[1][2] ), .C(n250), .D(\U2/x[0][2] ), .Q(
        \U2/n291 ) );
  INV3 U616 ( .A(\U2/n292 ), .Q(\U2/n13 ) );
  AOI221 U617 ( .A(n248), .B(\U2/x[1][1] ), .C(n262), .D(\U2/x[0][1] ), .Q(
        \U2/n292 ) );
  INV3 U618 ( .A(\U2/n293 ), .Q(\U2/n15 ) );
  AOI221 U619 ( .A(n245), .B(\U2/x[1][0] ), .C(n249), .D(\U2/x[0][0] ), .Q(
        \U2/n293 ) );
  INV3 U620 ( .A(\U2/n294 ), .Q(\U2/n17 ) );
  AOI221 U621 ( .A(n245), .B(\U2/x[2][7] ), .C(n262), .D(\U2/x[1][7] ), .Q(
        \U2/n294 ) );
  INV3 U622 ( .A(\U2/n295 ), .Q(\U2/n18 ) );
  AOI221 U623 ( .A(n245), .B(\U2/x[2][6] ), .C(n249), .D(\U2/x[1][6] ), .Q(
        \U2/n295 ) );
  INV3 U624 ( .A(\U2/n296 ), .Q(\U2/n19 ) );
  AOI221 U625 ( .A(n245), .B(\U2/x[2][5] ), .C(n250), .D(\U2/x[1][5] ), .Q(
        \U2/n296 ) );
  INV3 U626 ( .A(\U2/n297 ), .Q(\U2/n20 ) );
  AOI221 U627 ( .A(n245), .B(\U2/x[2][4] ), .C(n262), .D(\U2/x[1][4] ), .Q(
        \U2/n297 ) );
  INV3 U628 ( .A(\U2/n298 ), .Q(\U2/n21 ) );
  AOI221 U629 ( .A(n245), .B(\U2/x[2][3] ), .C(n262), .D(\U2/x[1][3] ), .Q(
        \U2/n298 ) );
  INV3 U630 ( .A(\U2/n299 ), .Q(\U2/n22 ) );
  AOI221 U631 ( .A(n245), .B(\U2/x[2][2] ), .C(n262), .D(\U2/x[1][2] ), .Q(
        \U2/n299 ) );
  INV3 U632 ( .A(\U2/n300 ), .Q(\U2/n23 ) );
  AOI221 U633 ( .A(n245), .B(\U2/x[2][1] ), .C(n261), .D(\U2/x[1][1] ), .Q(
        \U2/n300 ) );
  INV3 U634 ( .A(\U2/n301 ), .Q(\U2/n24 ) );
  AOI221 U635 ( .A(n245), .B(\U2/x[2][0] ), .C(n250), .D(\U2/x[1][0] ), .Q(
        \U2/n301 ) );
  INV3 U636 ( .A(\U2/n318 ), .Q(\U2/n226 ) );
  AOI221 U637 ( .A(n247), .B(\U2/x[28][7] ), .C(\U2/n286 ), .D(\U2/x[27][7] ), 
        .Q(\U2/n318 ) );
  INV3 U638 ( .A(\U2/n319 ), .Q(\U2/n228 ) );
  AOI221 U639 ( .A(n247), .B(\U2/x[28][6] ), .C(n250), .D(\U2/x[27][6] ), .Q(
        \U2/n319 ) );
  INV3 U640 ( .A(\U2/n320 ), .Q(\U2/n230 ) );
  AOI221 U641 ( .A(n247), .B(\U2/x[28][5] ), .C(n249), .D(\U2/x[27][5] ), .Q(
        \U2/n320 ) );
  INV3 U642 ( .A(\U2/n321 ), .Q(\U2/n232 ) );
  AOI221 U643 ( .A(\U2/n285 ), .B(\U2/x[28][4] ), .C(n261), .D(\U2/x[27][4] ), 
        .Q(\U2/n321 ) );
  INV3 U644 ( .A(\U2/n322 ), .Q(\U2/n234 ) );
  AOI221 U645 ( .A(\U2/n285 ), .B(\U2/x[28][3] ), .C(n249), .D(\U2/x[27][3] ), 
        .Q(\U2/n322 ) );
  INV3 U646 ( .A(\U2/n323 ), .Q(\U2/n236 ) );
  AOI221 U647 ( .A(\U2/n285 ), .B(\U2/x[28][2] ), .C(n262), .D(\U2/x[27][2] ), 
        .Q(\U2/n323 ) );
  INV3 U648 ( .A(\U2/n324 ), .Q(\U2/n238 ) );
  AOI221 U649 ( .A(n247), .B(\U2/x[28][1] ), .C(n249), .D(\U2/x[27][1] ), .Q(
        \U2/n324 ) );
  INV3 U650 ( .A(\U2/n325 ), .Q(\U2/n240 ) );
  AOI221 U651 ( .A(n247), .B(\U2/x[28][0] ), .C(n261), .D(\U2/x[27][0] ), .Q(
        \U2/n325 ) );
  INV3 U652 ( .A(\U2/n326 ), .Q(\U2/n241 ) );
  AOI221 U653 ( .A(\U2/n285 ), .B(\U2/x[29][7] ), .C(n249), .D(\U2/x[28][7] ), 
        .Q(\U2/n326 ) );
  INV3 U654 ( .A(\U2/n327 ), .Q(\U2/n242 ) );
  AOI221 U655 ( .A(n247), .B(\U2/x[29][6] ), .C(n249), .D(\U2/x[28][6] ), .Q(
        \U2/n327 ) );
  INV3 U656 ( .A(\U2/n328 ), .Q(\U2/n243 ) );
  AOI221 U657 ( .A(n248), .B(\U2/x[29][5] ), .C(n261), .D(\U2/x[28][5] ), .Q(
        \U2/n328 ) );
  INV3 U658 ( .A(\U2/n329 ), .Q(\U2/n244 ) );
  AOI221 U659 ( .A(n248), .B(\U2/x[29][4] ), .C(n261), .D(\U2/x[28][4] ), .Q(
        \U2/n329 ) );
  INV3 U660 ( .A(\U2/n330 ), .Q(\U2/n245 ) );
  AOI221 U661 ( .A(n245), .B(\U2/x[29][3] ), .C(\U2/n286 ), .D(\U2/x[28][3] ), 
        .Q(\U2/n330 ) );
  INV3 U662 ( .A(\U2/n331 ), .Q(\U2/n246 ) );
  AOI221 U663 ( .A(n247), .B(\U2/x[29][2] ), .C(n250), .D(\U2/x[28][2] ), .Q(
        \U2/n331 ) );
  INV3 U664 ( .A(\U2/n332 ), .Q(\U2/n247 ) );
  AOI221 U665 ( .A(n247), .B(\U2/x[29][1] ), .C(n261), .D(\U2/x[28][1] ), .Q(
        \U2/n332 ) );
  INV3 U666 ( .A(\U2/n333 ), .Q(\U2/n248 ) );
  AOI221 U667 ( .A(n247), .B(\U2/x[29][0] ), .C(n262), .D(\U2/x[28][0] ), .Q(
        \U2/n333 ) );
  INV3 U668 ( .A(\U2/n334 ), .Q(\U2/n249 ) );
  AOI221 U669 ( .A(n247), .B(\U2/x[30][7] ), .C(n249), .D(\U2/x[29][7] ), .Q(
        \U2/n334 ) );
  INV3 U670 ( .A(\U2/n335 ), .Q(\U2/n250 ) );
  AOI221 U671 ( .A(n248), .B(\U2/x[30][6] ), .C(n261), .D(\U2/x[29][6] ), .Q(
        \U2/n335 ) );
  INV3 U672 ( .A(\U2/n336 ), .Q(\U2/n251 ) );
  AOI221 U673 ( .A(n248), .B(\U2/x[30][5] ), .C(n262), .D(\U2/x[29][5] ), .Q(
        \U2/n336 ) );
  INV3 U674 ( .A(\U2/n337 ), .Q(\U2/n252 ) );
  AOI221 U675 ( .A(n248), .B(\U2/x[30][4] ), .C(n261), .D(\U2/x[29][4] ), .Q(
        \U2/n337 ) );
  INV3 U676 ( .A(\U2/n338 ), .Q(\U2/n253 ) );
  AOI221 U677 ( .A(n248), .B(\U2/x[30][3] ), .C(n261), .D(\U2/x[29][3] ), .Q(
        \U2/n338 ) );
  INV3 U678 ( .A(\U2/n339 ), .Q(\U2/n254 ) );
  AOI221 U679 ( .A(n248), .B(\U2/x[30][2] ), .C(n249), .D(\U2/x[29][2] ), .Q(
        \U2/n339 ) );
  INV3 U680 ( .A(\U2/n340 ), .Q(\U2/n255 ) );
  AOI221 U681 ( .A(n248), .B(\U2/x[30][1] ), .C(n250), .D(\U2/x[29][1] ), .Q(
        \U2/n340 ) );
  INV3 U682 ( .A(\U2/n341 ), .Q(\U2/n256 ) );
  AOI221 U683 ( .A(n248), .B(\U2/x[30][0] ), .C(n261), .D(\U2/x[29][0] ), .Q(
        \U2/n341 ) );
  INV3 U684 ( .A(\U2/n310 ), .Q(\U2/n257 ) );
  AOI221 U685 ( .A(n246), .B(\U2/x[31][7] ), .C(n262), .D(\U2/x[30][7] ), .Q(
        \U2/n310 ) );
  INV3 U686 ( .A(\U2/n311 ), .Q(\U2/n258 ) );
  AOI221 U687 ( .A(n246), .B(\U2/x[31][6] ), .C(n262), .D(\U2/x[30][6] ), .Q(
        \U2/n311 ) );
  INV3 U688 ( .A(\U2/n312 ), .Q(\U2/n259 ) );
  AOI221 U689 ( .A(n246), .B(\U2/x[31][5] ), .C(n262), .D(\U2/x[30][5] ), .Q(
        \U2/n312 ) );
  INV3 U690 ( .A(\U2/n313 ), .Q(\U2/n260 ) );
  AOI221 U691 ( .A(n246), .B(\U2/x[31][4] ), .C(n250), .D(\U2/x[30][4] ), .Q(
        \U2/n313 ) );
  INV3 U692 ( .A(\U2/n314 ), .Q(\U2/n261 ) );
  AOI221 U693 ( .A(n246), .B(\U2/x[31][3] ), .C(n250), .D(\U2/x[30][3] ), .Q(
        \U2/n314 ) );
  INV3 U694 ( .A(\U2/n315 ), .Q(\U2/n262 ) );
  AOI221 U695 ( .A(n247), .B(\U2/x[31][2] ), .C(n262), .D(\U2/x[30][2] ), .Q(
        \U2/n315 ) );
  INV3 U696 ( .A(\U2/n316 ), .Q(\U2/n263 ) );
  AOI221 U697 ( .A(n247), .B(\U2/x[31][1] ), .C(n262), .D(\U2/x[30][1] ), .Q(
        \U2/n316 ) );
  INV3 U698 ( .A(\U2/n317 ), .Q(\U2/n264 ) );
  AOI221 U699 ( .A(n247), .B(\U2/x[31][0] ), .C(n250), .D(\U2/x[30][0] ), .Q(
        \U2/n317 ) );
  NOR31 U700 ( .A(n121), .B(\U6/n33 ), .C(n19), .Q(\U6/n27 ) );
  NAND22 U701 ( .A(\U7/n9 ), .B(n148), .Q(\U7/n12 ) );
  NAND22 U702 ( .A(Filter_In[7]), .B(\U9/n3 ), .Q(\U9/n10 ) );
  NAND22 U703 ( .A(Filter_In[6]), .B(\U9/n3 ), .Q(\U9/n9 ) );
  NAND22 U704 ( .A(Filter_In[5]), .B(\U9/n3 ), .Q(\U9/n8 ) );
  NAND22 U705 ( .A(Filter_In[4]), .B(\U9/n3 ), .Q(\U9/n7 ) );
  NAND22 U706 ( .A(Filter_In[3]), .B(\U9/n3 ), .Q(\U9/n6 ) );
  NAND22 U707 ( .A(Filter_In[2]), .B(\U9/n3 ), .Q(\U9/n5 ) );
  NAND22 U708 ( .A(Filter_In[1]), .B(\U9/n3 ), .Q(\U9/n4 ) );
  NAND22 U709 ( .A(Filter_In[0]), .B(\U9/n3 ), .Q(\U9/n2 ) );
  NAND22 U710 ( .A(Accu_out[19]), .B(\U5/n3 ), .Q(\U5/n10 ) );
  NAND22 U711 ( .A(Accu_out[18]), .B(\U5/n3 ), .Q(\U5/n9 ) );
  NAND22 U712 ( .A(Accu_out[17]), .B(\U5/n3 ), .Q(\U5/n8 ) );
  NAND22 U713 ( .A(Accu_out[16]), .B(\U5/n3 ), .Q(\U5/n7 ) );
  NAND22 U714 ( .A(Accu_out[15]), .B(\U5/n3 ), .Q(\U5/n6 ) );
  NAND22 U715 ( .A(Accu_out[14]), .B(\U5/n3 ), .Q(\U5/n5 ) );
  NAND22 U716 ( .A(Accu_out[13]), .B(\U5/n3 ), .Q(\U5/n4 ) );
  NAND22 U717 ( .A(Accu_out[12]), .B(\U5/n3 ), .Q(\U5/n2 ) );
  NAND22 U718 ( .A(Accu_out[19]), .B(\U6/n24 ), .Q(
        \U4/mult_add_27_aco/PROD_not[19] ) );
  INV3 U719 ( .A(\U6/n25 ), .Q(\U6/n10 ) );
  AOI2111 U720 ( .A(\U6/n26 ), .B(\U6/n11 ), .C(Buff_OE), .D(ack_F2ADC), .Q(
        \U6/n25 ) );
  NAND31 U721 ( .A(\U6/n47 ), .B(\U6/n27 ), .C(\U6/n48 ), .Q(\U6/n26 ) );
  AOI211 U722 ( .A(n150), .B(\U7/n2 ), .C(n56), .Q(ADC_Rdb) );
  NOR31 U723 ( .A(n148), .B(\U7/n9 ), .C(n56), .Q(\U7/n13 ) );
  NOR31 U724 ( .A(\U8/n5 ), .B(\U8/pre_req_F2DAC ), .C(\U8/current_state ), 
        .Q(\U8/N5 ) );
  NOR21 U725 ( .A(n56), .B(\U7/n10 ), .Q(\U7/n15 ) );
  NOR21 U726 ( .A(ADC_Eocb), .B(n150), .Q(\U7/n11 ) );
  INV3 U727 ( .A(RESET), .Q(n263) );
  LOGIC0 U728 ( .Q(LDACb) );
  LOGIC1 U729 ( .Q(CLRb) );
endmodule

