/tp/xph2app/xph2app102/projet_Numerique/git/zigbee_project_2/implem/pnr/PNR_TOP_ANTHO_NETLIST_4/SCRIPTS/c35b4_A.lef