
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_FILTER is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_FILTER;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FILTER.all;

entity FILTER is

   port( Filter_In : in std_logic_vector (7 downto 0);  CLK, RESET, ADC_Eocb : 
         in std_logic;  ADC_Convstb, ADC_Rdb, ADC_csb, DAC_WRb, DAC_csb, LDACb,
         CLRb : out std_logic;  Filter_Out : out std_logic_vector (7 downto 0)
         );

end FILTER;

architecture SYN_A of FILTER is

   component LOGIC1
      port( Q : out std_logic);
   end component;
   
   component LOGIC0
      port( Q : out std_logic);
   end component;
   
   component INV3
      port( A : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR21
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR31
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI211
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND31
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI2111
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND22
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI221
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI2111
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND41
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component XNR21
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR22
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component BUF2
      port( A : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR40
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR21
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI311
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component IMUX21
      port( A, B, S : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND33
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI210
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND30
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND20
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI220
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR20
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component XNR20
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI220
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND21
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI211
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI221
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI310
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI210
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR20
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component INV2
      port( A : in std_logic;  Q : out std_logic);
   end component;
   
   component CLKIN3
      port( A : in std_logic;  Q : out std_logic);
   end component;
   
   component INV1
      port( A : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI222
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component CLKIN1
      port( A : in std_logic;  Q : out std_logic);
   end component;
   
   component IMAJ31
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI212
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component MUX22
      port( A, B, S : in std_logic;  Q : out std_logic);
   end component;
   
   component XNR31
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR30
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR31
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component ADD32
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DF3
      port( D, C : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFC3
      port( D, C, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal ADC_Rdb_port, DAC_WRb_port, Rom_Address_4_port, Rom_Address_3_port, 
      Rom_Address_2_port, Rom_Address_0_port, Rom_out_7_port, Rom_out_6_port, 
      Rom_out_5_port, Rom_out_4_port, Rom_out_3_port, Rom_out_2_port, 
      Rom_out_1_port, Rom_out_0_port, Filter_In_mem_7_port, 
      Filter_In_mem_6_port, Filter_In_mem_5_port, Filter_In_mem_4_port, 
      Filter_In_mem_3_port, Filter_In_mem_2_port, Filter_In_mem_1_port, 
      Filter_In_mem_0_port, Delay_Line_sample_shift, Delay_Line_out_6_port, 
      Delay_Line_out_3_port, Delay_Line_out_2_port, Delay_Line_out_1_port, 
      Mult_out_15_port, Mult_out_14_port, Mult_out_13_port, Mult_out_12_port, 
      Mult_out_11_port, Mult_out_10_port, Mult_out_9_port, Mult_out_8_port, 
      Mult_out_7_port, Mult_out_6_port, Mult_out_5_port, Mult_out_4_port, 
      Mult_out_3_port, Mult_out_2_port, Mult_out_1_port, Mult_out_0_port, 
      Accu_out_19_port, Accu_out_18_port, Accu_out_17_port, Accu_out_16_port, 
      Accu_out_15_port, Accu_out_14_port, Accu_out_13_port, Accu_out_12_port, 
      Buff_OE, req_ADC2F, ack_F2ADC, req_F2DAC, U1_n53, U1_n52, U1_n51, U1_n50,
      U1_n49, U1_n48, U1_n47, U1_n46, U1_n45, U1_n44, U1_n43, U1_n42, U1_n41, 
      U1_n40, U1_n39, U1_n38, U1_n37, U1_n36, U1_n35, U1_n34, U1_n33, U1_n32, 
      U1_n31, U1_n30, U1_n29, U1_n28, U1_n27, U1_n26, U1_n25, U1_n24, U1_n23, 
      U1_n22, U1_n21, U1_n20, U1_n19, U1_n18, U1_n17, U1_n16, U1_n15, U1_n14, 
      U1_n13, U1_n12, U1_n11, U1_n9, U1_n7, U1_n6, U1_n5, U1_n4, U1_n3, U1_n2, 
      U2_n741, U2_n740, U2_n739, U2_n738, U2_n737, U2_n736, U2_n735, U2_n734, 
      U2_n733, U2_n732, U2_n731, U2_n730, U2_n729, U2_n728, U2_n727, U2_n726, 
      U2_n725, U2_n724, U2_n723, U2_n722, U2_n721, U2_n720, U2_n719, U2_n718, 
      U2_n717, U2_n716, U2_n715, U2_n714, U2_n713, U2_n712, U2_n711, U2_n710, 
      U2_n709, U2_n708, U2_n707, U2_n706, U2_n705, U2_n704, U2_n703, U2_n702, 
      U2_n701, U2_n700, U2_n699, U2_n698, U2_n697, U2_n696, U2_n695, U2_n694, 
      U2_n693, U2_n692, U2_n691, U2_n690, U2_n689, U2_n688, U2_n687, U2_n686, 
      U2_n685, U2_n684, U2_n683, U2_n682, U2_n681, U2_n680, U2_n679, U2_n678, 
      U2_n677, U2_n676, U2_n675, U2_n674, U2_n673, U2_n672, U2_n671, U2_n670, 
      U2_n669, U2_n668, U2_n667, U2_n666, U2_n665, U2_n664, U2_n663, U2_n662, 
      U2_n661, U2_n660, U2_n659, U2_n658, U2_n657, U2_n656, U2_n655, U2_n654, 
      U2_n653, U2_n652, U2_n651, U2_n650, U2_n649, U2_n648, U2_n647, U2_n646, 
      U2_n645, U2_n644, U2_n643, U2_n642, U2_n641, U2_n640, U2_n639, U2_n638, 
      U2_n637, U2_n636, U2_n635, U2_n634, U2_n633, U2_n632, U2_n631, U2_n630, 
      U2_n629, U2_n628, U2_n627, U2_n626, U2_n625, U2_n624, U2_n623, U2_n622, 
      U2_n621, U2_n620, U2_n619, U2_n618, U2_n617, U2_n616, U2_n615, U2_n614, 
      U2_n613, U2_n612, U2_n611, U2_n610, U2_n609, U2_n608, U2_n607, U2_n606, 
      U2_n605, U2_n604, U2_n603, U2_n602, U2_n601, U2_n600, U2_n599, U2_n598, 
      U2_n597, U2_n596, U2_n595, U2_n594, U2_n593, U2_n592, U2_n523, U2_n522, 
      U2_n521, U2_n520, U2_n519, U2_n518, U2_n517, U2_n516, U2_n391, U2_n390, 
      U2_n389, U2_n388, U2_n387, U2_n386, U2_n385, U2_n384, U2_n383, U2_n382, 
      U2_n381, U2_n380, U2_n379, U2_n378, U2_n377, U2_n376, U2_n375, U2_n374, 
      U2_n373, U2_n372, U2_n371, U2_n370, U2_n369, U2_n368, U2_n367, U2_n366, 
      U2_n365, U2_n364, U2_n363, U2_n362, U2_n361, U2_n360, U2_n359, U2_n358, 
      U2_n357, U2_n356, U2_n355, U2_n354, U2_n353, U2_n352, U2_n351, U2_n350, 
      U2_n349, U2_n348, U2_n347, U2_n346, U2_n345, U2_n344, U2_n343, U2_n342, 
      U2_n341, U2_n340, U2_n339, U2_n338, U2_n337, U2_n336, U2_n335, U2_n334, 
      U2_n333, U2_n332, U2_n331, U2_n330, U2_n329, U2_n328, U2_n327, U2_n326, 
      U2_n325, U2_n324, U2_n323, U2_n322, U2_n321, U2_n320, U2_n319, U2_n318, 
      U2_n317, U2_n316, U2_n315, U2_n314, U2_n313, U2_n312, U2_n311, U2_n310, 
      U2_n309, U2_n308, U2_n307, U2_n306, U2_n305, U2_n304, U2_n303, U2_n302, 
      U2_n301, U2_n300, U2_n299, U2_n298, U2_n297, U2_n296, U2_n295, U2_n294, 
      U2_n293, U2_n292, U2_n291, U2_n290, U2_n289, U2_n288, U2_n287, U2_n286, 
      U2_n285, U2_n284, U2_n280, U2_n278, U2_n277, U2_n276, U2_n275, U2_n274, 
      U2_n273, U2_n272, U2_n271, U2_n270, U2_n269, U2_n268, U2_n267, U2_n266, 
      U2_n264, U2_n263, U2_n262, U2_n261, U2_n260, U2_n259, U2_n258, U2_n257, 
      U2_n256, U2_n255, U2_n254, U2_n253, U2_n252, U2_n251, U2_n250, U2_n249, 
      U2_n248, U2_n247, U2_n246, U2_n245, U2_n244, U2_n243, U2_n242, U2_n241, 
      U2_n240, U2_n238, U2_n236, U2_n234, U2_n232, U2_n230, U2_n228, U2_n226, 
      U2_n32, U2_n31, U2_n30, U2_n29, U2_n28, U2_n27, U2_n26, U2_n25, U2_n24, 
      U2_n23, U2_n22, U2_n21, U2_n20, U2_n19, U2_n18, U2_n17, U2_n16, U2_n15, 
      U2_n14, U2_n13, U2_n12, U2_n11, U2_n10, U2_n9, U2_n8, U2_n7, U2_n6, U2_n5
      , U2_n4, U2_n3, U2_n2, U2_n1, U2_n591, U2_n590, U2_n589, U2_n588, U2_n587
      , U2_n586, U2_n585, U2_n584, U2_n583, U2_n582, U2_n581, U2_n580, U2_n579,
      U2_n578, U2_n577, U2_n576, U2_n575, U2_n574, U2_n573, U2_n572, U2_n571, 
      U2_n570, U2_n569, U2_n568, U2_n567, U2_n566, U2_n565, U2_n564, U2_n563, 
      U2_n562, U2_n561, U2_n560, U2_n559, U2_n558, U2_n557, U2_n556, U2_n555, 
      U2_n554, U2_n553, U2_n552, U2_n551, U2_n550, U2_n549, U2_n548, U2_n547, 
      U2_n546, U2_n545, U2_n544, U2_n543, U2_n542, U2_n541, U2_n540, U2_n539, 
      U2_n538, U2_n537, U2_n536, U2_n535, U2_n534, U2_n533, U2_n532, U2_n531, 
      U2_n530, U2_n529, U2_n528, U2_n527, U2_n526, U2_n525, U2_n524, U2_n515, 
      U2_n514, U2_n513, U2_n512, U2_n511, U2_n510, U2_n509, U2_n508, U2_n507, 
      U2_n506, U2_n505, U2_n504, U2_n503, U2_n502, U2_n501, U2_n500, U2_n499, 
      U2_n498, U2_n497, U2_n496, U2_n495, U2_n494, U2_n493, U2_n492, U2_n491, 
      U2_n490, U2_n489, U2_n488, U2_n487, U2_n486, U2_n485, U2_n484, U2_n483, 
      U2_n482, U2_n481, U2_n480, U2_n479, U2_n478, U2_n477, U2_n476, U2_n475, 
      U2_n474, U2_n473, U2_n472, U2_n471, U2_n470, U2_n469, U2_n468, U2_n467, 
      U2_n466, U2_n465, U2_n464, U2_n463, U2_n462, U2_n461, U2_n460, U2_n459, 
      U2_n458, U2_n457, U2_n456, U2_n455, U2_n454, U2_n453, U2_n452, U2_n451, 
      U2_n450, U2_n449, U2_n448, U2_n447, U2_n446, U2_n445, U2_n444, U2_n443, 
      U2_n442, U2_n441, U2_n440, U2_n439, U2_n438, U2_n437, U2_n436, U2_n435, 
      U2_n434, U2_n433, U2_n432, U2_n431, U2_n430, U2_n429, U2_n428, U2_n427, 
      U2_n426, U2_n425, U2_n424, U2_n423, U2_n422, U2_n421, U2_n420, U2_n419, 
      U2_n418, U2_n417, U2_n416, U2_n415, U2_n414, U2_n413, U2_n412, U2_n411, 
      U2_n410, U2_n409, U2_n408, U2_n407, U2_n406, U2_n405, U2_n404, U2_n403, 
      U2_n402, U2_n401, U2_n400, U2_n399, U2_n398, U2_n397, U2_n396, U2_n395, 
      U2_n394, U2_n393, U2_n392, U2_x_31_0_port, U2_x_31_1_port, U2_x_31_2_port
      , U2_x_31_3_port, U2_x_31_4_port, U2_x_31_5_port, U2_x_31_6_port, 
      U2_x_31_7_port, U2_x_30_0_port, U2_x_30_1_port, U2_x_30_2_port, 
      U2_x_30_3_port, U2_x_30_4_port, U2_x_30_5_port, U2_x_30_6_port, 
      U2_x_30_7_port, U2_x_29_0_port, U2_x_29_1_port, U2_x_29_2_port, 
      U2_x_29_3_port, U2_x_29_4_port, U2_x_29_5_port, U2_x_29_6_port, 
      U2_x_29_7_port, U2_x_28_0_port, U2_x_28_1_port, U2_x_28_2_port, 
      U2_x_28_3_port, U2_x_28_4_port, U2_x_28_5_port, U2_x_28_6_port, 
      U2_x_28_7_port, U2_x_27_0_port, U2_x_27_1_port, U2_x_27_2_port, 
      U2_x_27_3_port, U2_x_27_4_port, U2_x_27_5_port, U2_x_27_6_port, 
      U2_x_27_7_port, U2_x_26_0_port, U2_x_26_1_port, U2_x_26_2_port, 
      U2_x_26_3_port, U2_x_26_4_port, U2_x_26_5_port, U2_x_26_6_port, 
      U2_x_26_7_port, U2_x_25_0_port, U2_x_25_1_port, U2_x_25_2_port, 
      U2_x_25_3_port, U2_x_25_4_port, U2_x_25_5_port, U2_x_25_6_port, 
      U2_x_25_7_port, U2_x_24_0_port, U2_x_24_1_port, U2_x_24_2_port, 
      U2_x_24_3_port, U2_x_24_4_port, U2_x_24_5_port, U2_x_24_6_port, 
      U2_x_24_7_port, U2_x_19_0_port, U2_x_19_1_port, U2_x_19_2_port, 
      U2_x_19_3_port, U2_x_19_4_port, U2_x_19_5_port, U2_x_19_6_port, 
      U2_x_19_7_port, U2_x_18_0_port, U2_x_18_1_port, U2_x_18_2_port, 
      U2_x_18_3_port, U2_x_18_4_port, U2_x_18_5_port, U2_x_18_6_port, 
      U2_x_18_7_port, U2_x_17_0_port, U2_x_17_1_port, U2_x_17_2_port, 
      U2_x_17_3_port, U2_x_17_4_port, U2_x_17_5_port, U2_x_17_6_port, 
      U2_x_17_7_port, U2_x_16_0_port, U2_x_16_1_port, U2_x_16_2_port, 
      U2_x_16_3_port, U2_x_16_4_port, U2_x_16_5_port, U2_x_16_6_port, 
      U2_x_16_7_port, U2_x_15_0_port, U2_x_15_1_port, U2_x_15_2_port, 
      U2_x_15_3_port, U2_x_15_4_port, U2_x_15_5_port, U2_x_15_6_port, 
      U2_x_15_7_port, U2_x_14_0_port, U2_x_14_1_port, U2_x_14_2_port, 
      U2_x_14_3_port, U2_x_14_4_port, U2_x_14_5_port, U2_x_14_6_port, 
      U2_x_14_7_port, U2_x_13_0_port, U2_x_13_1_port, U2_x_13_2_port, 
      U2_x_13_3_port, U2_x_13_4_port, U2_x_13_5_port, U2_x_13_6_port, 
      U2_x_13_7_port, U2_x_12_0_port, U2_x_12_1_port, U2_x_12_2_port, 
      U2_x_12_3_port, U2_x_12_4_port, U2_x_12_5_port, U2_x_12_6_port, 
      U2_x_12_7_port, U2_x_11_0_port, U2_x_11_1_port, U2_x_11_2_port, 
      U2_x_11_3_port, U2_x_11_4_port, U2_x_11_5_port, U2_x_11_6_port, 
      U2_x_11_7_port, U2_x_10_0_port, U2_x_10_1_port, U2_x_10_2_port, 
      U2_x_10_3_port, U2_x_10_4_port, U2_x_10_5_port, U2_x_10_6_port, 
      U2_x_10_7_port, U2_x_9_0_port, U2_x_9_1_port, U2_x_9_2_port, 
      U2_x_9_3_port, U2_x_9_4_port, U2_x_9_5_port, U2_x_9_6_port, U2_x_9_7_port
      , U2_x_8_0_port, U2_x_8_1_port, U2_x_8_2_port, U2_x_8_3_port, 
      U2_x_8_4_port, U2_x_8_5_port, U2_x_8_6_port, U2_x_8_7_port, U2_x_3_0_port
      , U2_x_3_1_port, U2_x_3_2_port, U2_x_3_3_port, U2_x_3_4_port, 
      U2_x_3_5_port, U2_x_3_6_port, U2_x_3_7_port, U2_x_2_0_port, U2_x_2_1_port
      , U2_x_2_2_port, U2_x_2_3_port, U2_x_2_4_port, U2_x_2_5_port, 
      U2_x_2_6_port, U2_x_2_7_port, U2_x_1_0_port, U2_x_1_1_port, U2_x_1_2_port
      , U2_x_1_3_port, U2_x_1_4_port, U2_x_1_5_port, U2_x_1_6_port, 
      U2_x_1_7_port, U2_x_0_0_port, U2_x_0_1_port, U2_x_0_2_port, U2_x_0_3_port
      , U2_x_0_4_port, U2_x_0_5_port, U2_x_0_6_port, U2_x_0_7_port, U4_n42, 
      U4_n41, U4_n40, U4_n39, U4_n38, U4_n37, U4_n36, U4_n35, U4_n34, U4_n33, 
      U4_n32, U4_n31, U4_n30, U4_n29, U4_n28, U4_N49, U4_N50, U4_N51, U4_N52, 
      U4_N53, U4_N54, U4_N55, U4_N56, U4_N57, U4_N58, U4_N59, U4_N60, U4_N61, 
      U4_N62, U4_N63, U4_N64, U4_N65, U4_N66, U4_N46, U4_N45, U4_N44, U4_N43, 
      U4_N42_port, U4_N41_port, U4_N40_port, U4_N39_port, U4_N38_port, 
      U4_N37_port, U4_N36_port, U4_N35_port, U4_N34_port, U4_N33_port, 
      U4_N32_port, U4_N31_port, U4_N30_port, U4_N29_port, U4_N28_port, U4_N27, 
      U4_N21, U4_N20, U4_N19, U4_N18, U4_N17, U4_N16, U4_N15, U4_N14, U4_N13, 
      U4_N12, U4_N11, U4_N10, U4_N9, U4_N8, U4_N7, U4_Accu_out_0_port, 
      U4_Accu_out_1_port, U4_Accu_out_2_port, U4_Accu_out_3_port, 
      U4_Accu_out_4_port, U4_Accu_out_5_port, U4_Accu_out_6_port, 
      U4_Accu_out_7_port, U4_Accu_out_8_port, U4_Accu_out_9_port, 
      U4_Accu_out_10_port, U4_Accu_out_11_port, U5_n11, U5_n10, U5_n9, U5_n8, 
      U5_n7, U5_n6, U5_n5, U5_n4, U5_n3, U5_n2, U5_n1, U5_n27, U5_n26, U5_n25, 
      U5_n24, U5_n23, U5_n22, U5_n21, U5_n20, U5_n19, U5_n18, U5_n17, U5_n16, 
      U5_n15, U5_n14, U5_n13, U5_n12, U6_n50, U6_n48, U6_n47, U6_n46, U6_n44, 
      U6_n43, U6_n36, U6_n35, U6_n34, U6_n32, U6_n31, U6_n29, U6_n28, U6_n27, 
      U6_n26, U6_n25, U6_n24, U6_n23, U6_n16, U6_n13, U6_n11, U6_n10, U6_n8, 
      U6_n7, U6_n33, U6_n4, U6_n2, U6_n42, U6_n41, U6_n40, U6_n39, U6_n38, 
      U6_n37, U6_n14, U7_n12, U7_n11, U7_n10, U7_n1, U7_n9, U7_n2, U7_n15, 
      U7_n14, U7_n13, U8_n5, U8_n1, U8_N5_port, U8_pre_req_F2DAC, 
      U8_current_state, U9_n11, U9_n10, U9_n9, U9_n8, U9_n7, U9_n6, U9_n5, 
      U9_n4, U9_n3, U9_n2, U9_n1, U9_n27, U9_n26, U9_n25, U9_n24, U9_n23, 
      U9_n22, U9_n21, U9_n20, U9_n19, U9_n18, U9_n17, U9_n16, U9_n15, U9_n14, 
      U9_n13, U9_n12, U3_mult_19_n91, U3_mult_19_n90, U3_mult_19_n89, 
      U3_mult_19_n88, U3_mult_19_n87, U3_mult_19_n86, U3_mult_19_n85, 
      U3_mult_19_n84, U3_mult_19_n83, U3_mult_19_n80, U3_mult_19_n79, 
      U3_mult_19_n78, U3_mult_19_n75, U3_mult_19_n72, U3_mult_19_n71, 
      U3_mult_19_n70, U3_mult_19_n67, U3_mult_19_n66, U3_mult_19_n65, 
      U3_mult_19_n64, U3_mult_19_n63, U3_mult_19_n62, U3_mult_19_n54, 
      U3_mult_19_n51, U3_mult_19_A2_7_port, U3_mult_19_A2_8_port, 
      U3_mult_19_A2_9_port, U3_mult_19_A2_10_port, U3_mult_19_A2_11_port, 
      U3_mult_19_A2_12_port, U3_mult_19_A1_7_port, U3_mult_19_A1_8_port, 
      U3_mult_19_A1_9_port, U3_mult_19_A1_10_port, U3_mult_19_A1_11_port, 
      U3_mult_19_A1_12_port, U3_mult_19_SUMB_1_1_port, U3_mult_19_SUMB_1_2_port
      , U3_mult_19_SUMB_1_3_port, U3_mult_19_SUMB_1_4_port, 
      U3_mult_19_SUMB_1_5_port, U3_mult_19_SUMB_1_6_port, 
      U3_mult_19_SUMB_2_1_port, U3_mult_19_SUMB_2_2_port, 
      U3_mult_19_SUMB_2_3_port, U3_mult_19_SUMB_2_4_port, 
      U3_mult_19_SUMB_2_5_port, U3_mult_19_SUMB_2_6_port, 
      U3_mult_19_SUMB_3_1_port, U3_mult_19_SUMB_3_2_port, 
      U3_mult_19_SUMB_3_3_port, U3_mult_19_SUMB_3_4_port, 
      U3_mult_19_SUMB_3_5_port, U3_mult_19_SUMB_3_6_port, 
      U3_mult_19_SUMB_4_1_port, U3_mult_19_SUMB_4_2_port, 
      U3_mult_19_SUMB_4_3_port, U3_mult_19_SUMB_4_4_port, 
      U3_mult_19_SUMB_4_5_port, U3_mult_19_SUMB_4_6_port, 
      U3_mult_19_SUMB_5_1_port, U3_mult_19_SUMB_5_2_port, 
      U3_mult_19_SUMB_5_3_port, U3_mult_19_SUMB_5_4_port, 
      U3_mult_19_SUMB_5_5_port, U3_mult_19_SUMB_5_6_port, 
      U3_mult_19_SUMB_6_1_port, U3_mult_19_SUMB_6_2_port, 
      U3_mult_19_SUMB_6_3_port, U3_mult_19_SUMB_6_4_port, 
      U3_mult_19_SUMB_6_5_port, U3_mult_19_SUMB_6_6_port, 
      U3_mult_19_SUMB_7_1_port, U3_mult_19_SUMB_7_2_port, 
      U3_mult_19_SUMB_7_3_port, U3_mult_19_SUMB_7_4_port, 
      U3_mult_19_SUMB_7_5_port, U3_mult_19_SUMB_7_6_port, 
      U3_mult_19_CARRYB_1_0_port, U3_mult_19_CARRYB_1_1_port, 
      U3_mult_19_CARRYB_1_2_port, U3_mult_19_CARRYB_1_3_port, 
      U3_mult_19_CARRYB_1_4_port, U3_mult_19_CARRYB_1_5_port, 
      U3_mult_19_CARRYB_1_6_port, U3_mult_19_CARRYB_2_0_port, 
      U3_mult_19_CARRYB_2_1_port, U3_mult_19_CARRYB_2_2_port, 
      U3_mult_19_CARRYB_2_3_port, U3_mult_19_CARRYB_2_4_port, 
      U3_mult_19_CARRYB_2_5_port, U3_mult_19_CARRYB_2_6_port, 
      U3_mult_19_CARRYB_3_0_port, U3_mult_19_CARRYB_3_1_port, 
      U3_mult_19_CARRYB_3_2_port, U3_mult_19_CARRYB_3_3_port, 
      U3_mult_19_CARRYB_3_4_port, U3_mult_19_CARRYB_3_5_port, 
      U3_mult_19_CARRYB_3_6_port, U3_mult_19_CARRYB_4_0_port, 
      U3_mult_19_CARRYB_4_1_port, U3_mult_19_CARRYB_4_2_port, 
      U3_mult_19_CARRYB_4_3_port, U3_mult_19_CARRYB_4_4_port, 
      U3_mult_19_CARRYB_4_5_port, U3_mult_19_CARRYB_4_6_port, 
      U3_mult_19_CARRYB_5_0_port, U3_mult_19_CARRYB_5_1_port, 
      U3_mult_19_CARRYB_5_2_port, U3_mult_19_CARRYB_5_3_port, 
      U3_mult_19_CARRYB_5_4_port, U3_mult_19_CARRYB_5_5_port, 
      U3_mult_19_CARRYB_5_6_port, U3_mult_19_CARRYB_6_0_port, 
      U3_mult_19_CARRYB_6_1_port, U3_mult_19_CARRYB_6_2_port, 
      U3_mult_19_CARRYB_6_3_port, U3_mult_19_CARRYB_6_4_port, 
      U3_mult_19_CARRYB_6_5_port, U3_mult_19_CARRYB_6_6_port, 
      U3_mult_19_CARRYB_7_0_port, U3_mult_19_CARRYB_7_1_port, 
      U3_mult_19_CARRYB_7_2_port, U3_mult_19_CARRYB_7_3_port, 
      U3_mult_19_CARRYB_7_4_port, U3_mult_19_CARRYB_7_5_port, 
      U3_mult_19_CARRYB_7_6_port, U3_mult_19_ab_0_1_port, 
      U3_mult_19_ab_0_2_port, U3_mult_19_ab_0_3_port, U3_mult_19_ab_0_4_port, 
      U3_mult_19_ab_0_5_port, U3_mult_19_ab_0_6_port, U3_mult_19_ab_0_7_port, 
      U3_mult_19_ab_1_0_port, U3_mult_19_ab_1_1_port, U3_mult_19_ab_1_2_port, 
      U3_mult_19_ab_1_3_port, U3_mult_19_ab_1_4_port, U3_mult_19_ab_1_5_port, 
      U3_mult_19_ab_1_6_port, U3_mult_19_ab_1_7_port, U3_mult_19_ab_2_0_port, 
      U3_mult_19_ab_2_1_port, U3_mult_19_ab_2_2_port, U3_mult_19_ab_2_3_port, 
      U3_mult_19_ab_2_4_port, U3_mult_19_ab_2_5_port, U3_mult_19_ab_2_6_port, 
      U3_mult_19_ab_2_7_port, U3_mult_19_ab_3_0_port, U3_mult_19_ab_3_1_port, 
      U3_mult_19_ab_3_2_port, U3_mult_19_ab_3_3_port, U3_mult_19_ab_3_4_port, 
      U3_mult_19_ab_3_5_port, U3_mult_19_ab_3_6_port, U3_mult_19_ab_3_7_port, 
      U3_mult_19_ab_4_0_port, U3_mult_19_ab_4_1_port, U3_mult_19_ab_4_2_port, 
      U3_mult_19_ab_4_3_port, U3_mult_19_ab_4_4_port, U3_mult_19_ab_4_5_port, 
      U3_mult_19_ab_4_6_port, U3_mult_19_ab_4_7_port, U3_mult_19_ab_5_0_port, 
      U3_mult_19_ab_5_1_port, U3_mult_19_ab_5_2_port, U3_mult_19_ab_5_3_port, 
      U3_mult_19_ab_5_4_port, U3_mult_19_ab_5_5_port, U3_mult_19_ab_5_6_port, 
      U3_mult_19_ab_5_7_port, U3_mult_19_ab_6_0_port, U3_mult_19_ab_6_1_port, 
      U3_mult_19_ab_6_2_port, U3_mult_19_ab_6_3_port, U3_mult_19_ab_6_4_port, 
      U3_mult_19_ab_6_5_port, U3_mult_19_ab_6_6_port, U3_mult_19_ab_6_7_port, 
      U3_mult_19_ab_7_0_port, U3_mult_19_ab_7_1_port, U3_mult_19_ab_7_2_port, 
      U3_mult_19_ab_7_3_port, U3_mult_19_ab_7_4_port, U3_mult_19_ab_7_5_port, 
      U3_mult_19_ab_7_6_port, U3_mult_19_ab_7_7_port, U4_add_27_aco_n20, 
      U4_add_27_aco_n18, U4_add_27_aco_n14, U4_add_27_aco_carry_1_port, 
      U4_add_27_aco_carry_2_port, U4_add_27_aco_carry_3_port, 
      U4_add_27_aco_carry_4_port, U4_add_27_aco_carry_5_port, 
      U4_add_27_aco_carry_6_port, U4_add_27_aco_carry_7_port, 
      U4_add_27_aco_carry_8_port, U4_add_27_aco_carry_9_port, 
      U4_add_27_aco_carry_10_port, U4_add_27_aco_carry_11_port, 
      U4_add_27_aco_carry_12_port, U4_add_27_aco_carry_13_port, 
      U4_add_27_aco_carry_14_port, U4_add_27_aco_carry_15_port, 
      U4_add_27_aco_carry_16_port, U4_add_27_aco_carry_17_port, 
      U4_add_27_aco_carry_18_port, U4_add_27_aco_carry_19_port, 
      U4_mult_add_27_aco_PROD_not_0_port, U4_mult_add_27_aco_PROD_not_1_port, 
      U4_mult_add_27_aco_PROD_not_2_port, U4_mult_add_27_aco_PROD_not_3_port, 
      U4_mult_add_27_aco_PROD_not_4_port, U4_mult_add_27_aco_PROD_not_5_port, 
      U4_mult_add_27_aco_PROD_not_6_port, U4_mult_add_27_aco_PROD_not_7_port, 
      U4_mult_add_27_aco_PROD_not_8_port, U4_mult_add_27_aco_PROD_not_9_port, 
      U4_mult_add_27_aco_PROD_not_10_port, U4_mult_add_27_aco_PROD_not_11_port,
      U4_mult_add_27_aco_PROD_not_12_port, U4_mult_add_27_aco_PROD_not_14_port,
      U4_mult_add_27_aco_PROD_not_15_port, U4_mult_add_27_aco_PROD_not_16_port,
      U4_mult_add_27_aco_PROD_not_17_port, U4_mult_add_27_aco_PROD_not_18_port,
      U4_mult_add_27_aco_PROD_not_19_port, U3_mult_19_FS_1_n39, 
      U3_mult_19_FS_1_n37, U3_mult_19_FS_1_n34, U3_mult_19_FS_1_n33, 
      U3_mult_19_FS_1_n32, U3_mult_19_FS_1_n31, U3_mult_19_FS_1_n29, 
      U3_mult_19_FS_1_n28, U3_mult_19_FS_1_n27, U3_mult_19_FS_1_n26, 
      U3_mult_19_FS_1_n25, U3_mult_19_FS_1_n24, U3_mult_19_FS_1_n23, 
      U3_mult_19_FS_1_n22, U3_mult_19_FS_1_n21, U3_mult_19_FS_1_n20, 
      U3_mult_19_FS_1_n19, U3_mult_19_FS_1_n18, U3_mult_19_FS_1_n17, 
      U3_mult_19_FS_1_n16, U3_mult_19_FS_1_n15, U3_mult_19_FS_1_n14, 
      U3_mult_19_FS_1_n13, U3_mult_19_FS_1_n12, U3_mult_19_FS_1_n11, 
      U3_mult_19_FS_1_n10, U3_mult_19_FS_1_n9, n3, n4, n5, n6, n7, n8, n9, n10,
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, 
      n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
      n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, 
      n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, 
      n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, 
      n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
      n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
      n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
      n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n_1000, 
      n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, 
      n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, 
      n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, 
      n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, 
      n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, 
      n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, 
      n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, 
      n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, 
      n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, 
      n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, 
      n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143 : 
      std_logic;

begin
   ADC_Rdb <= ADC_Rdb_port;
   ADC_csb <= ADC_Rdb_port;
   DAC_WRb <= DAC_WRb_port;
   DAC_csb <= DAC_WRb_port;
   
   U1_U27 : OAI212 port map( A => Rom_Address_4_port, B => U1_n48, C => U1_n49,
                           Q => Rom_out_1_port);
   U1_U26 : OAI212 port map( A => n232, B => U1_n29, C => U1_n7, Q => U1_n47);
   U1_U25 : OAI212 port map( A => n233, B => U1_n12, C => U1_n47, Q => U1_n44);
   U1_U14 : OAI222 port map( A => Rom_out_7_port, B => U1_n36, C => U1_n37, D 
                           => U1_n38, Q => Rom_out_3_port);
   U1_U7 : OAI212 port map( A => U1_n27, B => U1_n28, C => U1_n2, Q => U1_n21);
   U2_U413 : OAI222 port map( A => n123, B => U2_n358, C => n34, D => U2_n359, 
                           Q => U2_n692);
   U2_U412 : OAI222 port map( A => n122, B => U2_n356, C => n33, D => n235, Q 
                           => U2_n693);
   U2_U399 : OAI222 port map( A => Rom_Address_4_port, B => U2_n678, C => 
                           U2_n679, D => U1_n2, Q => Delay_Line_out_1_port);
   U2_U376 : OAI222 port map( A => Rom_Address_4_port, B => U2_n656, C => 
                           U2_n657, D => U1_n2, Q => Delay_Line_out_2_port);
   U2_U353 : OAI222 port map( A => Rom_Address_4_port, B => U2_n634, C => 
                           U2_n635, D => U1_n2, Q => Delay_Line_out_3_port);
   U2_U344 : OAI222 port map( A => n139, B => U2_n358, C => n51, D => n236, Q 
                           => U2_n626);
   U2_U343 : OAI222 port map( A => n138, B => U2_n356, C => n50, D => n235, Q 
                           => U2_n627);
   U2_U333 : OAI222 port map( A => n137, B => U2_n358, C => n49, D => n236, Q 
                           => U2_n616);
   U2_U332 : OAI222 port map( A => n25, B => U2_n356, C => n18, D => n235, Q =>
                           U2_n617);
   U2_U321 : OAI222 port map( A => n136, B => U2_n358, C => n48, D => n236, Q 
                           => U2_n604);
   U2_U320 : OAI222 port map( A => n135, B => U2_n356, C => n47, D => U2_n357, 
                           Q => U2_n605);
   U2_U310 : OAI222 port map( A => n134, B => U2_n358, C => n46, D => n236, Q 
                           => U2_n594);
   U2_U309 : OAI222 port map( A => n24, B => U2_n356, C => n17, D => U2_n357, Q
                           => U2_n595);
   U2_U298 : OAI222 port map( A => n147, B => U2_n358, C => n29, D => n236, Q 
                           => U2_n390);
   U2_U297 : OAI222 port map( A => n146, B => U2_n356, C => n55, D => U2_n357, 
                           Q => U2_n391);
   U2_U287 : OAI222 port map( A => n145, B => U2_n358, C => n54, D => n236, Q 
                           => U2_n380);
   U2_U286 : OAI222 port map( A => n144, B => U2_n356, C => n28, D => U2_n357, 
                           Q => U2_n381);
   U2_U284 : OAI222 port map( A => Rom_Address_4_port, B => U2_n376, C => 
                           U2_n377, D => U1_n2, Q => Delay_Line_out_6_port);
   U2_U275 : OAI222 port map( A => n143, B => U2_n358, C => n27, D => n236, Q 
                           => U2_n368);
   U2_U274 : OAI222 port map( A => n142, B => U2_n356, C => n53, D => U2_n357, 
                           Q => U2_n369);
   U2_U264 : OAI222 port map( A => n141, B => U2_n358, C => n52, D => n236, Q 
                           => U2_n354);
   U2_U263 : OAI222 port map( A => n140, B => U2_n356, C => n26, D => U2_n357, 
                           Q => U2_n355);
   U2_U226 : OAI222 port map( A => n238, B => n216, C => n251, D => n67, Q => 
                           U2_n392);
   U2_U225 : OAI222 port map( A => n239, B => n215, C => n251, D => n66, Q => 
                           U2_n393);
   U2_U224 : OAI222 port map( A => n240, B => n222, C => n251, D => n120, Q => 
                           U2_n394);
   U2_U223 : OAI222 port map( A => n239, B => n221, C => n251, D => n119, Q => 
                           U2_n395);
   U2_U222 : OAI222 port map( A => n240, B => n220, C => n251, D => n118, Q => 
                           U2_n396);
   U2_U221 : OAI222 port map( A => n241, B => n219, C => n251, D => n117, Q => 
                           U2_n397);
   U2_U220 : OAI222 port map( A => n244, B => n218, C => n252, D => n116, Q => 
                           U2_n398);
   U2_U219 : OAI222 port map( A => n244, B => n217, C => n252, D => n115, Q => 
                           U2_n399);
   U2_U218 : OAI222 port map( A => n241, B => n67, C => n252, D => n159, Q => 
                           U2_n400);
   U2_U217 : OAI222 port map( A => n242, B => n66, C => n252, D => n158, Q => 
                           U2_n401);
   U2_U216 : OAI222 port map( A => n241, B => n120, C => n252, D => n206, Q => 
                           U2_n402);
   U2_U215 : OAI222 port map( A => n242, B => n119, C => n252, D => n205, Q => 
                           U2_n403);
   U2_U214 : OAI222 port map( A => n244, B => n118, C => n253, D => n204, Q => 
                           U2_n404);
   U2_U213 : OAI222 port map( A => n244, B => n117, C => n253, D => n203, Q => 
                           U2_n405);
   U2_U212 : OAI222 port map( A => n243, B => n116, C => n253, D => n202, Q => 
                           U2_n406);
   U2_U211 : OAI222 port map( A => n240, B => n115, C => n253, D => n201, Q => 
                           U2_n407);
   U2_U210 : OAI222 port map( A => n237, B => n159, C => n253, D => n65, Q => 
                           U2_n408);
   U2_U209 : OAI222 port map( A => n238, B => n158, C => n253, D => n64, Q => 
                           U2_n409);
   U2_U208 : OAI222 port map( A => n240, B => n206, C => n254, D => n114, Q => 
                           U2_n410);
   U2_U207 : OAI222 port map( A => n238, B => n205, C => n254, D => n113, Q => 
                           U2_n411);
   U2_U206 : OAI222 port map( A => n240, B => n204, C => n254, D => n112, Q => 
                           U2_n412);
   U2_U205 : OAI222 port map( A => n241, B => n203, C => n254, D => n111, Q => 
                           U2_n413);
   U2_U204 : OAI222 port map( A => n242, B => n202, C => n254, D => n110, Q => 
                           U2_n414);
   U2_U203 : OAI222 port map( A => n242, B => n201, C => n254, D => n109, Q => 
                           U2_n415);
   U2_U202 : OAI222 port map( A => n243, B => n65, C => n251, D => n21, Q => 
                           U2_n416);
   U2_U201 : OAI222 port map( A => n243, B => n64, C => n252, D => n20, Q => 
                           U2_n417);
   U2_U200 : OAI222 port map( A => n244, B => n114, C => n253, D => n22, Q => 
                           U2_n418);
   U2_U199 : OAI222 port map( A => n244, B => n113, C => n254, D => n23, Q => 
                           U2_n419);
   U2_U198 : OAI222 port map( A => n244, B => n112, C => n253, D => n25, Q => 
                           U2_n420);
   U2_U197 : OAI222 port map( A => n243, B => n111, C => n254, D => n24, Q => 
                           U2_n421);
   U2_U196 : OAI222 port map( A => n242, B => n110, C => n255, D => n144, Q => 
                           U2_n422);
   U2_U195 : OAI222 port map( A => n242, B => n109, C => n255, D => n140, Q => 
                           U2_n423);
   U2_U194 : OAI222 port map( A => n241, B => n21, C => n255, D => n16, Q => 
                           U2_n424);
   U2_U193 : OAI222 port map( A => n243, B => n20, C => n255, D => n124, Q => 
                           U2_n425);
   U2_U192 : OAI222 port map( A => n239, B => n22, C => n255, D => n41, Q => 
                           U2_n426);
   U2_U191 : OAI222 port map( A => n240, B => n23, C => n255, D => n45, Q => 
                           U2_n427);
   U2_U190 : OAI222 port map( A => n243, B => n25, C => n253, D => n18, Q => 
                           U2_n428);
   U2_U189 : OAI222 port map( A => n244, B => n24, C => n252, D => n17, Q => 
                           U2_n429);
   U2_U188 : OAI222 port map( A => n240, B => n144, C => n255, D => n28, Q => 
                           U2_n430);
   U2_U187 : OAI222 port map( A => n237, B => n140, C => n256, D => n26, Q => 
                           U2_n431);
   U2_U186 : OAI222 port map( A => n242, B => n16, C => n255, D => n127, Q => 
                           U2_n432);
   U2_U185 : OAI222 port map( A => n238, B => n124, C => n256, D => n15, Q => 
                           U2_n433);
   U2_U184 : OAI222 port map( A => n241, B => n41, C => n256, D => n130, Q => 
                           U2_n434);
   U2_U183 : OAI222 port map( A => n240, B => n45, C => n256, D => n133, Q => 
                           U2_n435);
   U2_U182 : OAI222 port map( A => n242, B => n18, C => n256, D => n137, Q => 
                           U2_n436);
   U2_U181 : OAI222 port map( A => n239, B => n17, C => n256, D => n134, Q => 
                           U2_n437);
   U2_U180 : OAI222 port map( A => n241, B => n28, C => n256, D => n145, Q => 
                           U2_n438);
   U2_U179 : OAI222 port map( A => n237, B => n26, C => n256, D => n141, Q => 
                           U2_n439);
   U2_U178 : OAI222 port map( A => n242, B => n127, C => n251, D => n37, Q => 
                           U2_n440);
   U2_U177 : OAI222 port map( A => n241, B => n15, C => n252, D => n32, Q => 
                           U2_n441);
   U2_U176 : OAI222 port map( A => n244, B => n130, C => n257, D => n40, Q => 
                           U2_n442);
   U2_U175 : OAI222 port map( A => n241, B => n133, C => n258, D => n44, Q => 
                           U2_n443);
   U2_U174 : OAI222 port map( A => n242, B => n137, C => n257, D => n49, Q => 
                           U2_n444);
   U2_U173 : OAI222 port map( A => n243, B => n134, C => n258, D => n46, Q => 
                           U2_n445);
   U2_U172 : OAI222 port map( A => n244, B => n145, C => n257, D => n54, Q => 
                           U2_n446);
   U2_U171 : OAI222 port map( A => n243, B => n141, C => n257, D => n52, Q => 
                           U2_n447);
   U2_U170 : OAI222 port map( A => n243, B => n37, C => n257, D => n157, Q => 
                           U2_n448);
   U2_U169 : OAI222 port map( A => n239, B => n32, C => n257, D => n156, Q => 
                           U2_n449);
   U2_U168 : OAI222 port map( A => n240, B => n40, C => n257, D => n200, Q => 
                           U2_n450);
   U2_U167 : OAI222 port map( A => n241, B => n44, C => n257, D => n199, Q => 
                           U2_n451);
   U2_U166 : OAI222 port map( A => n244, B => n49, C => n258, D => n198, Q => 
                           U2_n452);
   U2_U165 : OAI222 port map( A => n239, B => n46, C => n258, D => n197, Q => 
                           U2_n453);
   U2_U164 : OAI222 port map( A => n238, B => n54, C => n258, D => n196, Q => 
                           U2_n454);
   U2_U163 : OAI222 port map( A => n242, B => n52, C => n258, D => n195, Q => 
                           U2_n455);
   U2_U162 : OAI222 port map( A => n243, B => n157, C => n258, D => n63, Q => 
                           U2_n456);
   U2_U161 : OAI222 port map( A => n243, B => n156, C => n258, D => n62, Q => 
                           U2_n457);
   U2_U160 : OAI222 port map( A => n241, B => n200, C => n255, D => n108, Q => 
                           U2_n458);
   U2_U159 : OAI222 port map( A => n238, B => n199, C => n251, D => n107, Q => 
                           U2_n459);
   U2_U158 : OAI222 port map( A => n239, B => n198, C => n259, D => n106, Q => 
                           U2_n460);
   U2_U157 : OAI222 port map( A => n240, B => n197, C => n254, D => n105, Q => 
                           U2_n461);
   U2_U156 : OAI222 port map( A => n238, B => n196, C => n259, D => n104, Q => 
                           U2_n462);
   U2_U155 : OAI222 port map( A => n239, B => n195, C => n259, D => n103, Q => 
                           U2_n463);
   U2_U154 : OAI222 port map( A => n238, B => n63, C => n259, D => n155, Q => 
                           U2_n464);
   U2_U153 : OAI222 port map( A => n244, B => n62, C => n259, D => n154, Q => 
                           U2_n465);
   U2_U152 : OAI222 port map( A => n244, B => n108, C => n259, D => n194, Q => 
                           U2_n466);
   U2_U151 : OAI222 port map( A => n238, B => n107, C => n259, D => n193, Q => 
                           U2_n467);
   U2_U150 : OAI222 port map( A => n241, B => n106, C => n259, D => n192, Q => 
                           U2_n468);
   U2_U149 : OAI222 port map( A => n239, B => n105, C => n259, D => n191, Q => 
                           U2_n469);
   U2_U148 : OAI222 port map( A => n243, B => n104, C => n259, D => n190, Q => 
                           U2_n470);
   U2_U147 : OAI222 port map( A => n244, B => n103, C => n251, D => n189, Q => 
                           U2_n471);
   U2_U146 : OAI222 port map( A => n237, B => n155, C => n259, D => n61, Q => 
                           U2_n472);
   U2_U145 : OAI222 port map( A => n237, B => n154, C => n258, D => n60, Q => 
                           U2_n473);
   U2_U144 : OAI222 port map( A => n237, B => n194, C => n252, D => n102, Q => 
                           U2_n474);
   U2_U143 : OAI222 port map( A => n237, B => n193, C => n253, D => n101, Q => 
                           U2_n475);
   U2_U142 : OAI222 port map( A => n237, B => n192, C => n260, D => n100, Q => 
                           U2_n476);
   U2_U141 : OAI222 port map( A => n238, B => n191, C => n251, D => n99, Q => 
                           U2_n477);
   U2_U140 : OAI222 port map( A => n238, B => n190, C => n252, D => n98, Q => 
                           U2_n478);
   U2_U139 : OAI222 port map( A => n238, B => n189, C => n259, D => n97, Q => 
                           U2_n479);
   U2_U138 : OAI222 port map( A => n238, B => n61, C => n254, D => n188, Q => 
                           U2_n480);
   U2_U137 : OAI222 port map( A => n238, B => n60, C => n251, D => n187, Q => 
                           U2_n481);
   U2_U136 : OAI222 port map( A => n237, B => n102, C => n254, D => n186, Q => 
                           U2_n482);
   U2_U135 : OAI222 port map( A => n237, B => n101, C => n257, D => n185, Q => 
                           U2_n483);
   U2_U134 : OAI222 port map( A => n238, B => n100, C => n258, D => n184, Q => 
                           U2_n484);
   U2_U133 : OAI222 port map( A => n239, B => n99, C => n259, D => n183, Q => 
                           U2_n485);
   U2_U132 : OAI222 port map( A => n240, B => n98, C => n260, D => n182, Q => 
                           U2_n486);
   U2_U131 : OAI222 port map( A => n238, B => n97, C => n257, D => n181, Q => 
                           U2_n487);
   U2_U130 : OAI222 port map( A => n237, B => n188, C => n255, D => n96, Q => 
                           U2_n488);
   U2_U129 : OAI222 port map( A => n238, B => n187, C => n256, D => n95, Q => 
                           U2_n489);
   U2_U128 : OAI222 port map( A => n239, B => n186, C => n257, D => n94, Q => 
                           U2_n490);
   U2_U127 : OAI222 port map( A => n240, B => n185, C => n258, D => n93, Q => 
                           U2_n491);
   U2_U126 : OAI222 port map( A => n239, B => n184, C => n253, D => n92, Q => 
                           U2_n492);
   U2_U125 : OAI222 port map( A => n239, B => n183, C => n254, D => n91, Q => 
                           U2_n493);
   U2_U124 : OAI222 port map( A => n239, B => n182, C => n258, D => n90, Q => 
                           U2_n494);
   U2_U123 : OAI222 port map( A => n239, B => n181, C => n253, D => n89, Q => 
                           U2_n495);
   U2_U122 : OAI222 port map( A => n239, B => n96, C => n254, D => n180, Q => 
                           U2_n496);
   U2_U121 : OAI222 port map( A => n240, B => n95, C => n251, D => n153, Q => 
                           U2_n497);
   U2_U120 : OAI222 port map( A => n240, B => n94, C => n252, D => n179, Q => 
                           U2_n498);
   U2_U119 : OAI222 port map( A => n240, B => n93, C => n255, D => n178, Q => 
                           U2_n499);
   U2_U118 : OAI222 port map( A => n240, B => n92, C => n252, D => n177, Q => 
                           U2_n500);
   U2_U117 : OAI222 port map( A => n240, B => n91, C => n255, D => n176, Q => 
                           U2_n501);
   U2_U116 : OAI222 port map( A => n238, B => n90, C => n256, D => n175, Q => 
                           U2_n502);
   U2_U115 : OAI222 port map( A => n241, B => n89, C => n257, D => n174, Q => 
                           U2_n503);
   U2_U114 : OAI222 port map( A => n238, B => n180, C => n258, D => n88, Q => 
                           U2_n504);
   U2_U113 : OAI222 port map( A => n242, B => n153, C => n253, D => n59, Q => 
                           U2_n505);
   U2_U112 : OAI222 port map( A => n242, B => n179, C => n260, D => n87, Q => 
                           U2_n506);
   U2_U111 : OAI222 port map( A => n237, B => n178, C => n260, D => n86, Q => 
                           U2_n507);
   U2_U110 : OAI222 port map( A => n239, B => n177, C => n260, D => n85, Q => 
                           U2_n508);
   U2_U109 : OAI222 port map( A => n244, B => n176, C => n260, D => n84, Q => 
                           U2_n509);
   U2_U108 : OAI222 port map( A => n244, B => n175, C => n260, D => n83, Q => 
                           U2_n510);
   U2_U107 : OAI222 port map( A => n237, B => n174, C => n260, D => n82, Q => 
                           U2_n511);
   U2_U106 : OAI222 port map( A => n243, B => n88, C => n257, D => n173, Q => 
                           U2_n512);
   U2_U105 : OAI222 port map( A => n243, B => n59, C => n259, D => n152, Q => 
                           U2_n513);
   U2_U104 : OAI222 port map( A => n238, B => n87, C => n258, D => n172, Q => 
                           U2_n514);
   U2_U103 : OAI222 port map( A => n237, B => n86, C => n259, D => n171, Q => 
                           U2_n515);
   U2_U94 : OAI222 port map( A => n238, B => n85, C => n251, D => n170, Q => 
                           U2_n524);
   U2_U93 : OAI222 port map( A => n244, B => n84, C => n253, D => n169, Q => 
                           U2_n525);
   U2_U92 : OAI222 port map( A => n239, B => n83, C => n254, D => n168, Q => 
                           U2_n526);
   U2_U91 : OAI222 port map( A => n243, B => n82, C => n257, D => n167, Q => 
                           U2_n527);
   U2_U90 : OAI222 port map( A => n240, B => n173, C => n258, D => n81, Q => 
                           U2_n528);
   U2_U89 : OAI222 port map( A => n240, B => n152, C => n252, D => n58, Q => 
                           U2_n529);
   U2_U88 : OAI222 port map( A => n242, B => n172, C => n253, D => n80, Q => 
                           U2_n530);
   U2_U87 : OAI222 port map( A => n240, B => n171, C => n258, D => n79, Q => 
                           U2_n531);
   U2_U86 : OAI222 port map( A => n243, B => n170, C => n253, D => n78, Q => 
                           U2_n532);
   U2_U85 : OAI222 port map( A => n242, B => n169, C => n253, D => n77, Q => 
                           U2_n533);
   U2_U84 : OAI222 port map( A => n238, B => n168, C => n253, D => n76, Q => 
                           U2_n534);
   U2_U83 : OAI222 port map( A => n240, B => n167, C => n254, D => n75, Q => 
                           U2_n535);
   U2_U82 : OAI222 port map( A => n242, B => n81, C => n259, D => n166, Q => 
                           U2_n536);
   U2_U81 : OAI222 port map( A => n237, B => n58, C => n254, D => n151, Q => 
                           U2_n537);
   U2_U80 : OAI222 port map( A => n238, B => n80, C => n260, D => n165, Q => 
                           U2_n538);
   U2_U79 : OAI222 port map( A => n241, B => n79, C => n260, D => n164, Q => 
                           U2_n539);
   U2_U78 : OAI222 port map( A => n241, B => n78, C => n253, D => n163, Q => 
                           U2_n540);
   U2_U77 : OAI222 port map( A => n241, B => n77, C => n260, D => n162, Q => 
                           U2_n541);
   U2_U76 : OAI222 port map( A => n241, B => n76, C => n252, D => n161, Q => 
                           U2_n542);
   U2_U75 : OAI222 port map( A => n241, B => n75, C => n258, D => n160, Q => 
                           U2_n543);
   U2_U74 : OAI222 port map( A => n241, B => n166, C => n255, D => n74, Q => 
                           U2_n544);
   U2_U73 : OAI222 port map( A => n242, B => n151, C => n254, D => n57, Q => 
                           U2_n545);
   U2_U72 : OAI222 port map( A => n242, B => n165, C => n260, D => n73, Q => 
                           U2_n546);
   U2_U71 : OAI222 port map( A => n242, B => n164, C => n255, D => n72, Q => 
                           U2_n547);
   U2_U70 : OAI222 port map( A => n242, B => n163, C => n256, D => n71, Q => 
                           U2_n548);
   U2_U69 : OAI222 port map( A => n242, B => n162, C => n260, D => n70, Q => 
                           U2_n549);
   U2_U68 : OAI222 port map( A => n243, B => n161, C => n256, D => n69, Q => 
                           U2_n550);
   U2_U67 : OAI222 port map( A => n243, B => n160, C => n257, D => n68, Q => 
                           U2_n551);
   U2_U66 : OAI222 port map( A => n243, B => n74, C => n258, D => n126, Q => 
                           U2_n552);
   U2_U65 : OAI222 port map( A => n243, B => n57, C => n259, D => n122, Q => 
                           U2_n553);
   U2_U64 : OAI222 port map( A => n243, B => n73, C => n256, D => n129, Q => 
                           U2_n554);
   U2_U63 : OAI222 port map( A => n239, B => n72, C => n255, D => n132, Q => 
                           U2_n555);
   U2_U62 : OAI222 port map( A => n239, B => n71, C => n255, D => n138, Q => 
                           U2_n556);
   U2_U61 : OAI222 port map( A => n237, B => n70, C => n256, D => n135, Q => 
                           U2_n557);
   U2_U60 : OAI222 port map( A => n238, B => n69, C => n260, D => n146, Q => 
                           U2_n558);
   U2_U59 : OAI222 port map( A => n237, B => n68, C => n256, D => n142, Q => 
                           U2_n559);
   U2_U58 : OAI222 port map( A => n244, B => n126, C => n256, D => n36, Q => 
                           U2_n560);
   U2_U57 : OAI222 port map( A => n244, B => n122, C => n259, D => n33, Q => 
                           U2_n561);
   U2_U56 : OAI222 port map( A => n244, B => n129, C => n251, D => n39, Q => 
                           U2_n562);
   U2_U55 : OAI222 port map( A => n244, B => n132, C => n251, D => n43, Q => 
                           U2_n563);
   U2_U54 : OAI222 port map( A => n244, B => n138, C => n256, D => n50, Q => 
                           U2_n564);
   U2_U53 : OAI222 port map( A => n237, B => n135, C => n254, D => n47, Q => 
                           U2_n565);
   U2_U52 : OAI222 port map( A => n243, B => n146, C => n260, D => n55, Q => 
                           U2_n566);
   U2_U51 : OAI222 port map( A => n237, B => n142, C => n252, D => n53, Q => 
                           U2_n567);
   U2_U50 : OAI222 port map( A => n241, B => n36, C => n252, D => n125, Q => 
                           U2_n568);
   U2_U49 : OAI222 port map( A => n242, B => n33, C => n251, D => n123, Q => 
                           U2_n569);
   U2_U48 : OAI222 port map( A => n239, B => n39, C => n251, D => n128, Q => 
                           U2_n570);
   U2_U47 : OAI222 port map( A => n240, B => n43, C => n257, D => n131, Q => 
                           U2_n571);
   U2_U46 : OAI222 port map( A => n237, B => n50, C => n254, D => n139, Q => 
                           U2_n572);
   U2_U45 : OAI222 port map( A => n237, B => n47, C => n257, D => n136, Q => 
                           U2_n573);
   U2_U44 : OAI222 port map( A => n239, B => n55, C => n255, D => n147, Q => 
                           U2_n574);
   U2_U43 : OAI222 port map( A => n242, B => n53, C => n256, D => n143, Q => 
                           U2_n575);
   U2_U42 : OAI222 port map( A => n244, B => n125, C => n257, D => n35, Q => 
                           U2_n576);
   U2_U41 : OAI222 port map( A => n241, B => n123, C => n258, D => n34, Q => 
                           U2_n577);
   U2_U40 : OAI222 port map( A => n242, B => n128, C => n259, D => n38, Q => 
                           U2_n578);
   U2_U39 : OAI222 port map( A => n244, B => n131, C => n251, D => n42, Q => 
                           U2_n579);
   U2_U38 : OAI222 port map( A => n239, B => n139, C => n260, D => n51, Q => 
                           U2_n580);
   U2_U37 : OAI222 port map( A => n240, B => n136, C => n254, D => n48, Q => 
                           U2_n581);
   U2_U36 : OAI222 port map( A => n241, B => n147, C => n259, D => n29, Q => 
                           U2_n582);
   U2_U35 : OAI222 port map( A => n237, B => n143, C => n260, D => n27, Q => 
                           U2_n583);
   U2_U34 : OAI222 port map( A => n243, B => n35, C => n253, D => n208, Q => 
                           U2_n584);
   U2_U33 : OAI222 port map( A => n239, B => n34, C => n252, D => n207, Q => 
                           U2_n585);
   U2_U32 : OAI222 port map( A => n237, B => n38, C => n252, D => n214, Q => 
                           U2_n586);
   U2_U31 : OAI222 port map( A => n240, B => n42, C => n260, D => n213, Q => 
                           U2_n587);
   U2_U30 : OAI222 port map( A => n241, B => n51, C => n255, D => n212, Q => 
                           U2_n588);
   U2_U29 : OAI222 port map( A => n241, B => n48, C => n260, D => n211, Q => 
                           U2_n589);
   U2_U28 : OAI222 port map( A => n243, B => n29, C => n257, D => n210, Q => 
                           U2_n590);
   U2_U27 : OAI222 port map( A => n237, B => n27, C => n260, D => n209, Q => 
                           U2_n591);
   U2_x_reg_31_0_inst : DF3 port map( D => U2_n264, C => CLK, Q => 
                           U2_x_31_0_port, QN => n_1000);
   U2_x_reg_31_1_inst : DF3 port map( D => U2_n263, C => CLK, Q => 
                           U2_x_31_1_port, QN => n_1001);
   U2_x_reg_31_2_inst : DF3 port map( D => U2_n262, C => CLK, Q => 
                           U2_x_31_2_port, QN => n_1002);
   U2_x_reg_31_3_inst : DF3 port map( D => U2_n261, C => CLK, Q => 
                           U2_x_31_3_port, QN => n_1003);
   U2_x_reg_31_4_inst : DF3 port map( D => U2_n260, C => CLK, Q => 
                           U2_x_31_4_port, QN => n_1004);
   U2_x_reg_31_5_inst : DF3 port map( D => U2_n259, C => CLK, Q => 
                           U2_x_31_5_port, QN => n_1005);
   U2_x_reg_31_6_inst : DF3 port map( D => U2_n258, C => CLK, Q => 
                           U2_x_31_6_port, QN => n_1006);
   U2_x_reg_31_7_inst : DF3 port map( D => U2_n257, C => CLK, Q => 
                           U2_x_31_7_port, QN => n_1007);
   U2_x_reg_30_0_inst : DF3 port map( D => U2_n256, C => CLK, Q => 
                           U2_x_30_0_port, QN => n_1008);
   U2_x_reg_30_1_inst : DF3 port map( D => U2_n255, C => CLK, Q => 
                           U2_x_30_1_port, QN => n_1009);
   U2_x_reg_30_2_inst : DF3 port map( D => U2_n254, C => CLK, Q => 
                           U2_x_30_2_port, QN => n_1010);
   U2_x_reg_30_3_inst : DF3 port map( D => U2_n253, C => CLK, Q => 
                           U2_x_30_3_port, QN => n_1011);
   U2_x_reg_30_4_inst : DF3 port map( D => U2_n252, C => CLK, Q => 
                           U2_x_30_4_port, QN => n_1012);
   U2_x_reg_30_5_inst : DF3 port map( D => U2_n251, C => CLK, Q => 
                           U2_x_30_5_port, QN => n_1013);
   U2_x_reg_30_6_inst : DF3 port map( D => U2_n250, C => CLK, Q => 
                           U2_x_30_6_port, QN => n_1014);
   U2_x_reg_30_7_inst : DF3 port map( D => U2_n249, C => CLK, Q => 
                           U2_x_30_7_port, QN => n_1015);
   U2_x_reg_29_0_inst : DF3 port map( D => U2_n248, C => CLK, Q => 
                           U2_x_29_0_port, QN => n_1016);
   U2_x_reg_29_1_inst : DF3 port map( D => U2_n247, C => CLK, Q => 
                           U2_x_29_1_port, QN => n_1017);
   U2_x_reg_29_2_inst : DF3 port map( D => U2_n246, C => CLK, Q => 
                           U2_x_29_2_port, QN => n_1018);
   U2_x_reg_29_3_inst : DF3 port map( D => U2_n245, C => CLK, Q => 
                           U2_x_29_3_port, QN => n_1019);
   U2_x_reg_29_4_inst : DF3 port map( D => U2_n244, C => CLK, Q => 
                           U2_x_29_4_port, QN => n_1020);
   U2_x_reg_29_5_inst : DF3 port map( D => U2_n243, C => CLK, Q => 
                           U2_x_29_5_port, QN => n_1021);
   U2_x_reg_29_6_inst : DF3 port map( D => U2_n242, C => CLK, Q => 
                           U2_x_29_6_port, QN => n_1022);
   U2_x_reg_29_7_inst : DF3 port map( D => U2_n241, C => CLK, Q => 
                           U2_x_29_7_port, QN => n_1023);
   U2_x_reg_28_0_inst : DF3 port map( D => U2_n240, C => CLK, Q => 
                           U2_x_28_0_port, QN => n_1024);
   U2_x_reg_28_1_inst : DF3 port map( D => U2_n238, C => CLK, Q => 
                           U2_x_28_1_port, QN => n_1025);
   U2_x_reg_28_2_inst : DF3 port map( D => U2_n236, C => CLK, Q => 
                           U2_x_28_2_port, QN => n_1026);
   U2_x_reg_28_3_inst : DF3 port map( D => U2_n234, C => CLK, Q => 
                           U2_x_28_3_port, QN => n_1027);
   U2_x_reg_28_4_inst : DF3 port map( D => U2_n232, C => CLK, Q => 
                           U2_x_28_4_port, QN => n_1028);
   U2_x_reg_28_5_inst : DF3 port map( D => U2_n230, C => CLK, Q => 
                           U2_x_28_5_port, QN => n_1029);
   U2_x_reg_28_6_inst : DF3 port map( D => U2_n228, C => CLK, Q => 
                           U2_x_28_6_port, QN => n_1030);
   U2_x_reg_28_7_inst : DF3 port map( D => U2_n226, C => CLK, Q => 
                           U2_x_28_7_port, QN => n_1031);
   U2_x_reg_27_0_inst : DF3 port map( D => U2_n392, C => CLK, Q => 
                           U2_x_27_0_port, QN => n216);
   U2_x_reg_27_1_inst : DF3 port map( D => U2_n393, C => CLK, Q => 
                           U2_x_27_1_port, QN => n215);
   U2_x_reg_27_2_inst : DF3 port map( D => U2_n394, C => CLK, Q => 
                           U2_x_27_2_port, QN => n222);
   U2_x_reg_27_3_inst : DF3 port map( D => U2_n395, C => CLK, Q => 
                           U2_x_27_3_port, QN => n221);
   U2_x_reg_27_4_inst : DF3 port map( D => U2_n396, C => CLK, Q => 
                           U2_x_27_4_port, QN => n220);
   U2_x_reg_27_5_inst : DF3 port map( D => U2_n397, C => CLK, Q => 
                           U2_x_27_5_port, QN => n219);
   U2_x_reg_27_6_inst : DF3 port map( D => U2_n398, C => CLK, Q => 
                           U2_x_27_6_port, QN => n218);
   U2_x_reg_27_7_inst : DF3 port map( D => U2_n399, C => CLK, Q => 
                           U2_x_27_7_port, QN => n217);
   U2_x_reg_26_0_inst : DF3 port map( D => U2_n400, C => CLK, Q => 
                           U2_x_26_0_port, QN => n67);
   U2_x_reg_26_1_inst : DF3 port map( D => U2_n401, C => CLK, Q => 
                           U2_x_26_1_port, QN => n66);
   U2_x_reg_26_2_inst : DF3 port map( D => U2_n402, C => CLK, Q => 
                           U2_x_26_2_port, QN => n120);
   U2_x_reg_26_3_inst : DF3 port map( D => U2_n403, C => CLK, Q => 
                           U2_x_26_3_port, QN => n119);
   U2_x_reg_26_4_inst : DF3 port map( D => U2_n404, C => CLK, Q => 
                           U2_x_26_4_port, QN => n118);
   U2_x_reg_26_5_inst : DF3 port map( D => U2_n405, C => CLK, Q => 
                           U2_x_26_5_port, QN => n117);
   U2_x_reg_26_6_inst : DF3 port map( D => U2_n406, C => CLK, Q => 
                           U2_x_26_6_port, QN => n116);
   U2_x_reg_26_7_inst : DF3 port map( D => U2_n407, C => CLK, Q => 
                           U2_x_26_7_port, QN => n115);
   U2_x_reg_25_0_inst : DF3 port map( D => U2_n408, C => CLK, Q => 
                           U2_x_25_0_port, QN => n159);
   U2_x_reg_25_1_inst : DF3 port map( D => U2_n409, C => CLK, Q => 
                           U2_x_25_1_port, QN => n158);
   U2_x_reg_25_2_inst : DF3 port map( D => U2_n410, C => CLK, Q => 
                           U2_x_25_2_port, QN => n206);
   U2_x_reg_25_3_inst : DF3 port map( D => U2_n411, C => CLK, Q => 
                           U2_x_25_3_port, QN => n205);
   U2_x_reg_25_4_inst : DF3 port map( D => U2_n412, C => CLK, Q => 
                           U2_x_25_4_port, QN => n204);
   U2_x_reg_25_5_inst : DF3 port map( D => U2_n413, C => CLK, Q => 
                           U2_x_25_5_port, QN => n203);
   U2_x_reg_25_6_inst : DF3 port map( D => U2_n414, C => CLK, Q => 
                           U2_x_25_6_port, QN => n202);
   U2_x_reg_25_7_inst : DF3 port map( D => U2_n415, C => CLK, Q => 
                           U2_x_25_7_port, QN => n201);
   U2_x_reg_24_0_inst : DF3 port map( D => U2_n416, C => CLK, Q => 
                           U2_x_24_0_port, QN => n65);
   U2_x_reg_24_1_inst : DF3 port map( D => U2_n417, C => CLK, Q => 
                           U2_x_24_1_port, QN => n64);
   U2_x_reg_24_2_inst : DF3 port map( D => U2_n418, C => CLK, Q => 
                           U2_x_24_2_port, QN => n114);
   U2_x_reg_24_3_inst : DF3 port map( D => U2_n419, C => CLK, Q => 
                           U2_x_24_3_port, QN => n113);
   U2_x_reg_24_4_inst : DF3 port map( D => U2_n420, C => CLK, Q => 
                           U2_x_24_4_port, QN => n112);
   U2_x_reg_24_5_inst : DF3 port map( D => U2_n421, C => CLK, Q => 
                           U2_x_24_5_port, QN => n111);
   U2_x_reg_24_6_inst : DF3 port map( D => U2_n422, C => CLK, Q => 
                           U2_x_24_6_port, QN => n110);
   U2_x_reg_24_7_inst : DF3 port map( D => U2_n423, C => CLK, Q => 
                           U2_x_24_7_port, QN => n109);
   U2_x_reg_23_0_inst : DF3 port map( D => U2_n424, C => CLK, Q => n_1032, QN 
                           => n21);
   U2_x_reg_23_1_inst : DF3 port map( D => U2_n425, C => CLK, Q => n_1033, QN 
                           => n20);
   U2_x_reg_23_2_inst : DF3 port map( D => U2_n426, C => CLK, Q => n_1034, QN 
                           => n22);
   U2_x_reg_23_3_inst : DF3 port map( D => U2_n427, C => CLK, Q => n_1035, QN 
                           => n23);
   U2_x_reg_23_4_inst : DF3 port map( D => U2_n428, C => CLK, Q => n_1036, QN 
                           => n25);
   U2_x_reg_23_5_inst : DF3 port map( D => U2_n429, C => CLK, Q => n_1037, QN 
                           => n24);
   U2_x_reg_23_6_inst : DF3 port map( D => U2_n430, C => CLK, Q => n_1038, QN 
                           => n144);
   U2_x_reg_23_7_inst : DF3 port map( D => U2_n431, C => CLK, Q => n_1039, QN 
                           => n140);
   U2_x_reg_22_0_inst : DF3 port map( D => U2_n432, C => CLK, Q => n_1040, QN 
                           => n16);
   U2_x_reg_22_1_inst : DF3 port map( D => U2_n433, C => CLK, Q => n_1041, QN 
                           => n124);
   U2_x_reg_22_2_inst : DF3 port map( D => U2_n434, C => CLK, Q => n_1042, QN 
                           => n41);
   U2_x_reg_22_3_inst : DF3 port map( D => U2_n435, C => CLK, Q => n_1043, QN 
                           => n45);
   U2_x_reg_22_4_inst : DF3 port map( D => U2_n436, C => CLK, Q => n_1044, QN 
                           => n18);
   U2_x_reg_22_5_inst : DF3 port map( D => U2_n437, C => CLK, Q => n_1045, QN 
                           => n17);
   U2_x_reg_22_6_inst : DF3 port map( D => U2_n438, C => CLK, Q => n_1046, QN 
                           => n28);
   U2_x_reg_22_7_inst : DF3 port map( D => U2_n439, C => CLK, Q => n_1047, QN 
                           => n26);
   U2_x_reg_21_0_inst : DF3 port map( D => U2_n440, C => CLK, Q => n_1048, QN 
                           => n127);
   U2_x_reg_21_1_inst : DF3 port map( D => U2_n441, C => CLK, Q => n_1049, QN 
                           => n15);
   U2_x_reg_21_2_inst : DF3 port map( D => U2_n442, C => CLK, Q => n_1050, QN 
                           => n130);
   U2_x_reg_21_3_inst : DF3 port map( D => U2_n443, C => CLK, Q => n_1051, QN 
                           => n133);
   U2_x_reg_21_4_inst : DF3 port map( D => U2_n444, C => CLK, Q => n_1052, QN 
                           => n137);
   U2_x_reg_21_5_inst : DF3 port map( D => U2_n445, C => CLK, Q => n_1053, QN 
                           => n134);
   U2_x_reg_21_6_inst : DF3 port map( D => U2_n446, C => CLK, Q => n_1054, QN 
                           => n145);
   U2_x_reg_21_7_inst : DF3 port map( D => U2_n447, C => CLK, Q => n_1055, QN 
                           => n141);
   U2_x_reg_20_0_inst : DF3 port map( D => U2_n448, C => CLK, Q => n_1056, QN 
                           => n37);
   U2_x_reg_20_1_inst : DF3 port map( D => U2_n449, C => CLK, Q => n_1057, QN 
                           => n32);
   U2_x_reg_20_2_inst : DF3 port map( D => U2_n450, C => CLK, Q => n_1058, QN 
                           => n40);
   U2_x_reg_20_3_inst : DF3 port map( D => U2_n451, C => CLK, Q => n_1059, QN 
                           => n44);
   U2_x_reg_20_4_inst : DF3 port map( D => U2_n452, C => CLK, Q => n_1060, QN 
                           => n49);
   U2_x_reg_20_5_inst : DF3 port map( D => U2_n453, C => CLK, Q => n_1061, QN 
                           => n46);
   U2_x_reg_20_6_inst : DF3 port map( D => U2_n454, C => CLK, Q => n_1062, QN 
                           => n54);
   U2_x_reg_20_7_inst : DF3 port map( D => U2_n455, C => CLK, Q => n_1063, QN 
                           => n52);
   U2_x_reg_19_0_inst : DF3 port map( D => U2_n456, C => CLK, Q => 
                           U2_x_19_0_port, QN => n157);
   U2_x_reg_19_1_inst : DF3 port map( D => U2_n457, C => CLK, Q => 
                           U2_x_19_1_port, QN => n156);
   U2_x_reg_19_2_inst : DF3 port map( D => U2_n458, C => CLK, Q => 
                           U2_x_19_2_port, QN => n200);
   U2_x_reg_19_3_inst : DF3 port map( D => U2_n459, C => CLK, Q => 
                           U2_x_19_3_port, QN => n199);
   U2_x_reg_19_4_inst : DF3 port map( D => U2_n460, C => CLK, Q => 
                           U2_x_19_4_port, QN => n198);
   U2_x_reg_19_5_inst : DF3 port map( D => U2_n461, C => CLK, Q => 
                           U2_x_19_5_port, QN => n197);
   U2_x_reg_19_6_inst : DF3 port map( D => U2_n462, C => CLK, Q => 
                           U2_x_19_6_port, QN => n196);
   U2_x_reg_19_7_inst : DF3 port map( D => U2_n463, C => CLK, Q => 
                           U2_x_19_7_port, QN => n195);
   U2_x_reg_18_0_inst : DF3 port map( D => U2_n464, C => CLK, Q => 
                           U2_x_18_0_port, QN => n63);
   U2_x_reg_18_1_inst : DF3 port map( D => U2_n465, C => CLK, Q => 
                           U2_x_18_1_port, QN => n62);
   U2_x_reg_18_2_inst : DF3 port map( D => U2_n466, C => CLK, Q => 
                           U2_x_18_2_port, QN => n108);
   U2_x_reg_18_3_inst : DF3 port map( D => U2_n467, C => CLK, Q => 
                           U2_x_18_3_port, QN => n107);
   U2_x_reg_18_4_inst : DF3 port map( D => U2_n468, C => CLK, Q => 
                           U2_x_18_4_port, QN => n106);
   U2_x_reg_18_5_inst : DF3 port map( D => U2_n469, C => CLK, Q => 
                           U2_x_18_5_port, QN => n105);
   U2_x_reg_18_6_inst : DF3 port map( D => U2_n470, C => CLK, Q => 
                           U2_x_18_6_port, QN => n104);
   U2_x_reg_18_7_inst : DF3 port map( D => U2_n471, C => CLK, Q => 
                           U2_x_18_7_port, QN => n103);
   U2_x_reg_17_0_inst : DF3 port map( D => U2_n472, C => CLK, Q => 
                           U2_x_17_0_port, QN => n155);
   U2_x_reg_17_1_inst : DF3 port map( D => U2_n473, C => CLK, Q => 
                           U2_x_17_1_port, QN => n154);
   U2_x_reg_17_2_inst : DF3 port map( D => U2_n474, C => CLK, Q => 
                           U2_x_17_2_port, QN => n194);
   U2_x_reg_17_3_inst : DF3 port map( D => U2_n475, C => CLK, Q => 
                           U2_x_17_3_port, QN => n193);
   U2_x_reg_17_4_inst : DF3 port map( D => U2_n476, C => CLK, Q => 
                           U2_x_17_4_port, QN => n192);
   U2_x_reg_17_5_inst : DF3 port map( D => U2_n477, C => CLK, Q => 
                           U2_x_17_5_port, QN => n191);
   U2_x_reg_17_6_inst : DF3 port map( D => U2_n478, C => CLK, Q => 
                           U2_x_17_6_port, QN => n190);
   U2_x_reg_17_7_inst : DF3 port map( D => U2_n479, C => CLK, Q => 
                           U2_x_17_7_port, QN => n189);
   U2_x_reg_16_0_inst : DF3 port map( D => U2_n480, C => CLK, Q => 
                           U2_x_16_0_port, QN => n61);
   U2_x_reg_16_1_inst : DF3 port map( D => U2_n481, C => CLK, Q => 
                           U2_x_16_1_port, QN => n60);
   U2_x_reg_16_2_inst : DF3 port map( D => U2_n482, C => CLK, Q => 
                           U2_x_16_2_port, QN => n102);
   U2_x_reg_16_3_inst : DF3 port map( D => U2_n483, C => CLK, Q => 
                           U2_x_16_3_port, QN => n101);
   U2_x_reg_16_4_inst : DF3 port map( D => U2_n484, C => CLK, Q => 
                           U2_x_16_4_port, QN => n100);
   U2_x_reg_16_5_inst : DF3 port map( D => U2_n485, C => CLK, Q => 
                           U2_x_16_5_port, QN => n99);
   U2_x_reg_16_6_inst : DF3 port map( D => U2_n486, C => CLK, Q => 
                           U2_x_16_6_port, QN => n98);
   U2_x_reg_16_7_inst : DF3 port map( D => U2_n487, C => CLK, Q => 
                           U2_x_16_7_port, QN => n97);
   U2_x_reg_15_0_inst : DF3 port map( D => U2_n488, C => CLK, Q => 
                           U2_x_15_0_port, QN => n188);
   U2_x_reg_15_1_inst : DF3 port map( D => U2_n489, C => CLK, Q => 
                           U2_x_15_1_port, QN => n187);
   U2_x_reg_15_2_inst : DF3 port map( D => U2_n490, C => CLK, Q => 
                           U2_x_15_2_port, QN => n186);
   U2_x_reg_15_3_inst : DF3 port map( D => U2_n491, C => CLK, Q => 
                           U2_x_15_3_port, QN => n185);
   U2_x_reg_15_4_inst : DF3 port map( D => U2_n492, C => CLK, Q => 
                           U2_x_15_4_port, QN => n184);
   U2_x_reg_15_5_inst : DF3 port map( D => U2_n493, C => CLK, Q => 
                           U2_x_15_5_port, QN => n183);
   U2_x_reg_15_6_inst : DF3 port map( D => U2_n494, C => CLK, Q => 
                           U2_x_15_6_port, QN => n182);
   U2_x_reg_15_7_inst : DF3 port map( D => U2_n495, C => CLK, Q => 
                           U2_x_15_7_port, QN => n181);
   U2_x_reg_14_0_inst : DF3 port map( D => U2_n496, C => CLK, Q => 
                           U2_x_14_0_port, QN => n96);
   U2_x_reg_14_1_inst : DF3 port map( D => U2_n497, C => CLK, Q => 
                           U2_x_14_1_port, QN => n95);
   U2_x_reg_14_2_inst : DF3 port map( D => U2_n498, C => CLK, Q => 
                           U2_x_14_2_port, QN => n94);
   U2_x_reg_14_3_inst : DF3 port map( D => U2_n499, C => CLK, Q => 
                           U2_x_14_3_port, QN => n93);
   U2_x_reg_14_4_inst : DF3 port map( D => U2_n500, C => CLK, Q => 
                           U2_x_14_4_port, QN => n92);
   U2_x_reg_14_5_inst : DF3 port map( D => U2_n501, C => CLK, Q => 
                           U2_x_14_5_port, QN => n91);
   U2_x_reg_14_6_inst : DF3 port map( D => U2_n502, C => CLK, Q => 
                           U2_x_14_6_port, QN => n90);
   U2_x_reg_14_7_inst : DF3 port map( D => U2_n503, C => CLK, Q => 
                           U2_x_14_7_port, QN => n89);
   U2_x_reg_13_0_inst : DF3 port map( D => U2_n504, C => CLK, Q => 
                           U2_x_13_0_port, QN => n180);
   U2_x_reg_13_1_inst : DF3 port map( D => U2_n505, C => CLK, Q => 
                           U2_x_13_1_port, QN => n153);
   U2_x_reg_13_2_inst : DF3 port map( D => U2_n506, C => CLK, Q => 
                           U2_x_13_2_port, QN => n179);
   U2_x_reg_13_3_inst : DF3 port map( D => U2_n507, C => CLK, Q => 
                           U2_x_13_3_port, QN => n178);
   U2_x_reg_13_4_inst : DF3 port map( D => U2_n508, C => CLK, Q => 
                           U2_x_13_4_port, QN => n177);
   U2_x_reg_13_5_inst : DF3 port map( D => U2_n509, C => CLK, Q => 
                           U2_x_13_5_port, QN => n176);
   U2_x_reg_13_6_inst : DF3 port map( D => U2_n510, C => CLK, Q => 
                           U2_x_13_6_port, QN => n175);
   U2_x_reg_13_7_inst : DF3 port map( D => U2_n511, C => CLK, Q => 
                           U2_x_13_7_port, QN => n174);
   U2_x_reg_12_0_inst : DF3 port map( D => U2_n512, C => CLK, Q => 
                           U2_x_12_0_port, QN => n88);
   U2_x_reg_12_1_inst : DF3 port map( D => U2_n513, C => CLK, Q => 
                           U2_x_12_1_port, QN => n59);
   U2_x_reg_12_2_inst : DF3 port map( D => U2_n514, C => CLK, Q => 
                           U2_x_12_2_port, QN => n87);
   U2_x_reg_12_3_inst : DF3 port map( D => U2_n515, C => CLK, Q => 
                           U2_x_12_3_port, QN => n86);
   U2_x_reg_12_4_inst : DF3 port map( D => U2_n524, C => CLK, Q => 
                           U2_x_12_4_port, QN => n85);
   U2_x_reg_12_5_inst : DF3 port map( D => U2_n525, C => CLK, Q => 
                           U2_x_12_5_port, QN => n84);
   U2_x_reg_12_6_inst : DF3 port map( D => U2_n526, C => CLK, Q => 
                           U2_x_12_6_port, QN => n83);
   U2_x_reg_12_7_inst : DF3 port map( D => U2_n527, C => CLK, Q => 
                           U2_x_12_7_port, QN => n82);
   U2_x_reg_11_0_inst : DF3 port map( D => U2_n528, C => CLK, Q => 
                           U2_x_11_0_port, QN => n173);
   U2_x_reg_11_1_inst : DF3 port map( D => U2_n529, C => CLK, Q => 
                           U2_x_11_1_port, QN => n152);
   U2_x_reg_11_2_inst : DF3 port map( D => U2_n530, C => CLK, Q => 
                           U2_x_11_2_port, QN => n172);
   U2_x_reg_11_3_inst : DF3 port map( D => U2_n531, C => CLK, Q => 
                           U2_x_11_3_port, QN => n171);
   U2_x_reg_11_4_inst : DF3 port map( D => U2_n532, C => CLK, Q => 
                           U2_x_11_4_port, QN => n170);
   U2_x_reg_11_5_inst : DF3 port map( D => U2_n533, C => CLK, Q => 
                           U2_x_11_5_port, QN => n169);
   U2_x_reg_11_6_inst : DF3 port map( D => U2_n534, C => CLK, Q => 
                           U2_x_11_6_port, QN => n168);
   U2_x_reg_11_7_inst : DF3 port map( D => U2_n535, C => CLK, Q => 
                           U2_x_11_7_port, QN => n167);
   U2_x_reg_10_0_inst : DF3 port map( D => U2_n536, C => CLK, Q => 
                           U2_x_10_0_port, QN => n81);
   U2_x_reg_10_1_inst : DF3 port map( D => U2_n537, C => CLK, Q => 
                           U2_x_10_1_port, QN => n58);
   U2_x_reg_10_2_inst : DF3 port map( D => U2_n538, C => CLK, Q => 
                           U2_x_10_2_port, QN => n80);
   U2_x_reg_10_3_inst : DF3 port map( D => U2_n539, C => CLK, Q => 
                           U2_x_10_3_port, QN => n79);
   U2_x_reg_10_4_inst : DF3 port map( D => U2_n540, C => CLK, Q => 
                           U2_x_10_4_port, QN => n78);
   U2_x_reg_10_5_inst : DF3 port map( D => U2_n541, C => CLK, Q => 
                           U2_x_10_5_port, QN => n77);
   U2_x_reg_10_6_inst : DF3 port map( D => U2_n542, C => CLK, Q => 
                           U2_x_10_6_port, QN => n76);
   U2_x_reg_10_7_inst : DF3 port map( D => U2_n543, C => CLK, Q => 
                           U2_x_10_7_port, QN => n75);
   U2_x_reg_9_0_inst : DF3 port map( D => U2_n544, C => CLK, Q => U2_x_9_0_port
                           , QN => n166);
   U2_x_reg_9_1_inst : DF3 port map( D => U2_n545, C => CLK, Q => U2_x_9_1_port
                           , QN => n151);
   U2_x_reg_9_2_inst : DF3 port map( D => U2_n546, C => CLK, Q => U2_x_9_2_port
                           , QN => n165);
   U2_x_reg_9_3_inst : DF3 port map( D => U2_n547, C => CLK, Q => U2_x_9_3_port
                           , QN => n164);
   U2_x_reg_9_4_inst : DF3 port map( D => U2_n548, C => CLK, Q => U2_x_9_4_port
                           , QN => n163);
   U2_x_reg_9_5_inst : DF3 port map( D => U2_n549, C => CLK, Q => U2_x_9_5_port
                           , QN => n162);
   U2_x_reg_9_6_inst : DF3 port map( D => U2_n550, C => CLK, Q => U2_x_9_6_port
                           , QN => n161);
   U2_x_reg_9_7_inst : DF3 port map( D => U2_n551, C => CLK, Q => U2_x_9_7_port
                           , QN => n160);
   U2_x_reg_8_0_inst : DF3 port map( D => U2_n552, C => CLK, Q => U2_x_8_0_port
                           , QN => n74);
   U2_x_reg_8_1_inst : DF3 port map( D => U2_n553, C => CLK, Q => U2_x_8_1_port
                           , QN => n57);
   U2_x_reg_8_2_inst : DF3 port map( D => U2_n554, C => CLK, Q => U2_x_8_2_port
                           , QN => n73);
   U2_x_reg_8_3_inst : DF3 port map( D => U2_n555, C => CLK, Q => U2_x_8_3_port
                           , QN => n72);
   U2_x_reg_8_4_inst : DF3 port map( D => U2_n556, C => CLK, Q => U2_x_8_4_port
                           , QN => n71);
   U2_x_reg_8_5_inst : DF3 port map( D => U2_n557, C => CLK, Q => U2_x_8_5_port
                           , QN => n70);
   U2_x_reg_8_6_inst : DF3 port map( D => U2_n558, C => CLK, Q => U2_x_8_6_port
                           , QN => n69);
   U2_x_reg_8_7_inst : DF3 port map( D => U2_n559, C => CLK, Q => U2_x_8_7_port
                           , QN => n68);
   U2_x_reg_7_0_inst : DF3 port map( D => U2_n560, C => CLK, Q => n_1064, QN =>
                           n126);
   U2_x_reg_7_1_inst : DF3 port map( D => U2_n561, C => CLK, Q => n_1065, QN =>
                           n122);
   U2_x_reg_7_2_inst : DF3 port map( D => U2_n562, C => CLK, Q => n_1066, QN =>
                           n129);
   U2_x_reg_7_3_inst : DF3 port map( D => U2_n563, C => CLK, Q => n_1067, QN =>
                           n132);
   U2_x_reg_7_4_inst : DF3 port map( D => U2_n564, C => CLK, Q => n_1068, QN =>
                           n138);
   U2_x_reg_7_5_inst : DF3 port map( D => U2_n565, C => CLK, Q => n_1069, QN =>
                           n135);
   U2_x_reg_7_6_inst : DF3 port map( D => U2_n566, C => CLK, Q => n_1070, QN =>
                           n146);
   U2_x_reg_7_7_inst : DF3 port map( D => U2_n567, C => CLK, Q => n_1071, QN =>
                           n142);
   U2_x_reg_6_0_inst : DF3 port map( D => U2_n568, C => CLK, Q => n_1072, QN =>
                           n36);
   U2_x_reg_6_1_inst : DF3 port map( D => U2_n569, C => CLK, Q => n_1073, QN =>
                           n33);
   U2_x_reg_6_2_inst : DF3 port map( D => U2_n570, C => CLK, Q => n_1074, QN =>
                           n39);
   U2_x_reg_6_3_inst : DF3 port map( D => U2_n571, C => CLK, Q => n_1075, QN =>
                           n43);
   U2_x_reg_6_4_inst : DF3 port map( D => U2_n572, C => CLK, Q => n_1076, QN =>
                           n50);
   U2_x_reg_6_5_inst : DF3 port map( D => U2_n573, C => CLK, Q => n_1077, QN =>
                           n47);
   U2_x_reg_6_6_inst : DF3 port map( D => U2_n574, C => CLK, Q => n_1078, QN =>
                           n55);
   U2_x_reg_6_7_inst : DF3 port map( D => U2_n575, C => CLK, Q => n_1079, QN =>
                           n53);
   U2_x_reg_5_0_inst : DF3 port map( D => U2_n576, C => CLK, Q => n_1080, QN =>
                           n125);
   U2_x_reg_5_1_inst : DF3 port map( D => U2_n577, C => CLK, Q => n_1081, QN =>
                           n123);
   U2_x_reg_5_2_inst : DF3 port map( D => U2_n578, C => CLK, Q => n_1082, QN =>
                           n128);
   U2_x_reg_5_3_inst : DF3 port map( D => U2_n579, C => CLK, Q => n_1083, QN =>
                           n131);
   U2_x_reg_5_4_inst : DF3 port map( D => U2_n580, C => CLK, Q => n_1084, QN =>
                           n139);
   U2_x_reg_5_5_inst : DF3 port map( D => U2_n581, C => CLK, Q => n_1085, QN =>
                           n136);
   U2_x_reg_5_6_inst : DF3 port map( D => U2_n582, C => CLK, Q => n_1086, QN =>
                           n147);
   U2_x_reg_5_7_inst : DF3 port map( D => U2_n583, C => CLK, Q => n_1087, QN =>
                           n143);
   U2_x_reg_4_0_inst : DF3 port map( D => U2_n584, C => CLK, Q => n_1088, QN =>
                           n35);
   U2_x_reg_4_1_inst : DF3 port map( D => U2_n585, C => CLK, Q => n_1089, QN =>
                           n34);
   U2_x_reg_4_2_inst : DF3 port map( D => U2_n586, C => CLK, Q => n_1090, QN =>
                           n38);
   U2_x_reg_4_3_inst : DF3 port map( D => U2_n587, C => CLK, Q => n_1091, QN =>
                           n42);
   U2_x_reg_4_4_inst : DF3 port map( D => U2_n588, C => CLK, Q => n_1092, QN =>
                           n51);
   U2_x_reg_4_5_inst : DF3 port map( D => U2_n589, C => CLK, Q => n_1093, QN =>
                           n48);
   U2_x_reg_4_6_inst : DF3 port map( D => U2_n590, C => CLK, Q => n_1094, QN =>
                           n29);
   U2_x_reg_4_7_inst : DF3 port map( D => U2_n591, C => CLK, Q => n_1095, QN =>
                           n27);
   U2_x_reg_3_0_inst : DF3 port map( D => U2_n32, C => CLK, Q => U2_x_3_0_port,
                           QN => n208);
   U2_x_reg_3_1_inst : DF3 port map( D => U2_n31, C => CLK, Q => U2_x_3_1_port,
                           QN => n207);
   U2_x_reg_3_2_inst : DF3 port map( D => U2_n30, C => CLK, Q => U2_x_3_2_port,
                           QN => n214);
   U2_x_reg_3_3_inst : DF3 port map( D => U2_n29, C => CLK, Q => U2_x_3_3_port,
                           QN => n213);
   U2_x_reg_3_4_inst : DF3 port map( D => U2_n28, C => CLK, Q => U2_x_3_4_port,
                           QN => n212);
   U2_x_reg_3_5_inst : DF3 port map( D => U2_n27, C => CLK, Q => U2_x_3_5_port,
                           QN => n211);
   U2_x_reg_3_6_inst : DF3 port map( D => U2_n26, C => CLK, Q => U2_x_3_6_port,
                           QN => n210);
   U2_x_reg_3_7_inst : DF3 port map( D => U2_n25, C => CLK, Q => U2_x_3_7_port,
                           QN => n209);
   U2_x_reg_2_0_inst : DF3 port map( D => U2_n24, C => CLK, Q => U2_x_2_0_port,
                           QN => n_1096);
   U2_x_reg_2_1_inst : DF3 port map( D => U2_n23, C => CLK, Q => U2_x_2_1_port,
                           QN => n_1097);
   U2_x_reg_2_2_inst : DF3 port map( D => U2_n22, C => CLK, Q => U2_x_2_2_port,
                           QN => n_1098);
   U2_x_reg_2_3_inst : DF3 port map( D => U2_n21, C => CLK, Q => U2_x_2_3_port,
                           QN => n_1099);
   U2_x_reg_2_4_inst : DF3 port map( D => U2_n20, C => CLK, Q => U2_x_2_4_port,
                           QN => n_1100);
   U2_x_reg_2_5_inst : DF3 port map( D => U2_n19, C => CLK, Q => U2_x_2_5_port,
                           QN => n_1101);
   U2_x_reg_2_6_inst : DF3 port map( D => U2_n18, C => CLK, Q => U2_x_2_6_port,
                           QN => n_1102);
   U2_x_reg_2_7_inst : DF3 port map( D => U2_n17, C => CLK, Q => U2_x_2_7_port,
                           QN => n_1103);
   U2_x_reg_1_0_inst : DF3 port map( D => U2_n15, C => CLK, Q => U2_x_1_0_port,
                           QN => n_1104);
   U2_x_reg_1_1_inst : DF3 port map( D => U2_n13, C => CLK, Q => U2_x_1_1_port,
                           QN => n_1105);
   U2_x_reg_1_2_inst : DF3 port map( D => U2_n11, C => CLK, Q => U2_x_1_2_port,
                           QN => n_1106);
   U2_x_reg_1_3_inst : DF3 port map( D => U2_n9, C => CLK, Q => U2_x_1_3_port, 
                           QN => n_1107);
   U2_x_reg_1_4_inst : DF3 port map( D => U2_n7, C => CLK, Q => U2_x_1_4_port, 
                           QN => n_1108);
   U2_x_reg_1_5_inst : DF3 port map( D => U2_n5, C => CLK, Q => U2_x_1_5_port, 
                           QN => n_1109);
   U2_x_reg_1_6_inst : DF3 port map( D => U2_n3, C => CLK, Q => U2_x_1_6_port, 
                           QN => n_1110);
   U2_x_reg_1_7_inst : DF3 port map( D => U2_n1, C => CLK, Q => U2_x_1_7_port, 
                           QN => n_1111);
   U2_x_reg_0_0_inst : DF3 port map( D => U2_n16, C => CLK, Q => U2_x_0_0_port,
                           QN => n_1112);
   U2_x_reg_0_1_inst : DF3 port map( D => U2_n14, C => CLK, Q => U2_x_0_1_port,
                           QN => n_1113);
   U2_x_reg_0_2_inst : DF3 port map( D => U2_n12, C => CLK, Q => U2_x_0_2_port,
                           QN => n_1114);
   U2_x_reg_0_3_inst : DF3 port map( D => U2_n10, C => CLK, Q => U2_x_0_3_port,
                           QN => n_1115);
   U2_x_reg_0_4_inst : DF3 port map( D => U2_n8, C => CLK, Q => U2_x_0_4_port, 
                           QN => n_1116);
   U2_x_reg_0_5_inst : DF3 port map( D => U2_n6, C => CLK, Q => U2_x_0_5_port, 
                           QN => n_1117);
   U2_x_reg_0_6_inst : DF3 port map( D => U2_n4, C => CLK, Q => U2_x_0_6_port, 
                           QN => n_1118);
   U2_x_reg_0_7_inst : DF3 port map( D => U2_n2, C => CLK, Q => U2_x_0_7_port, 
                           QN => n_1119);
   U4_ACCU_reg_19_inst : DF3 port map( D => U4_N46, C => CLK, Q => 
                           Accu_out_19_port, QN => n_1120);
   U4_ACCU_reg_18_inst : DF3 port map( D => U4_N45, C => CLK, Q => 
                           Accu_out_18_port, QN => n_1121);
   U4_ACCU_reg_17_inst : DF3 port map( D => U4_N44, C => CLK, Q => 
                           Accu_out_17_port, QN => n_1122);
   U4_ACCU_reg_16_inst : DF3 port map( D => U4_N43, C => CLK, Q => 
                           Accu_out_16_port, QN => n_1123);
   U4_ACCU_reg_15_inst : DF3 port map( D => U4_N42_port, C => CLK, Q => 
                           Accu_out_15_port, QN => n_1124);
   U4_ACCU_reg_14_inst : DF3 port map( D => U4_N41_port, C => CLK, Q => 
                           Accu_out_14_port, QN => n_1125);
   U4_ACCU_reg_13_inst : DF3 port map( D => U4_N40_port, C => CLK, Q => 
                           Accu_out_13_port, QN => n8);
   U4_ACCU_reg_12_inst : DF3 port map( D => U4_N39_port, C => CLK, Q => 
                           Accu_out_12_port, QN => n_1126);
   U4_ACCU_reg_11_inst : DF3 port map( D => U4_N38_port, C => CLK, Q => 
                           U4_Accu_out_11_port, QN => n_1127);
   U4_ACCU_reg_10_inst : DF3 port map( D => U4_N37_port, C => CLK, Q => 
                           U4_Accu_out_10_port, QN => n_1128);
   U4_ACCU_reg_9_inst : DF3 port map( D => U4_N36_port, C => CLK, Q => 
                           U4_Accu_out_9_port, QN => n_1129);
   U4_ACCU_reg_8_inst : DF3 port map( D => U4_N35_port, C => CLK, Q => 
                           U4_Accu_out_8_port, QN => n_1130);
   U4_ACCU_reg_7_inst : DF3 port map( D => U4_N34_port, C => CLK, Q => 
                           U4_Accu_out_7_port, QN => n_1131);
   U4_ACCU_reg_6_inst : DF3 port map( D => U4_N33_port, C => CLK, Q => 
                           U4_Accu_out_6_port, QN => n_1132);
   U4_ACCU_reg_5_inst : DF3 port map( D => U4_N32_port, C => CLK, Q => 
                           U4_Accu_out_5_port, QN => n_1133);
   U4_ACCU_reg_4_inst : DF3 port map( D => U4_N31_port, C => CLK, Q => 
                           U4_Accu_out_4_port, QN => n_1134);
   U4_ACCU_reg_3_inst : DF3 port map( D => U4_N30_port, C => CLK, Q => 
                           U4_Accu_out_3_port, QN => n_1135);
   U4_ACCU_reg_2_inst : DF3 port map( D => U4_N29_port, C => CLK, Q => 
                           U4_Accu_out_2_port, QN => n_1136);
   U4_ACCU_reg_1_inst : DF3 port map( D => U4_N28_port, C => CLK, Q => 
                           U4_Accu_out_1_port, QN => n_1137);
   U4_ACCU_reg_0_inst : DF3 port map( D => U4_N27, C => CLK, Q => 
                           U4_Accu_out_0_port, QN => n_1138);
   U5_U17 : OAI212 port map( A => U5_n19, B => U5_n1, C => U5_n10, Q => U5_n20)
                           ;
   U5_U15 : OAI212 port map( A => U5_n18, B => U5_n1, C => U5_n9, Q => U5_n21);
   U5_U13 : OAI212 port map( A => U5_n17, B => U5_n1, C => U5_n8, Q => U5_n22);
   U5_U11 : OAI212 port map( A => U5_n16, B => U5_n1, C => U5_n7, Q => U5_n23);
   U5_U9 : OAI212 port map( A => U5_n15, B => U5_n1, C => U5_n6, Q => U5_n24);
   U5_U7 : OAI212 port map( A => U5_n14, B => U5_n1, C => U5_n5, Q => U5_n25);
   U5_U5 : OAI212 port map( A => U5_n13, B => U5_n1, C => U5_n4, Q => U5_n26);
   U5_U3 : OAI212 port map( A => U5_n12, B => U5_n1, C => U5_n2, Q => U5_n27);
   U5_Buff_out_reg_0_inst : DF3 port map( D => U5_n27, C => CLK, Q => 
                           Filter_Out(0), QN => U5_n12);
   U5_Buff_out_reg_1_inst : DF3 port map( D => U5_n26, C => CLK, Q => 
                           Filter_Out(1), QN => U5_n13);
   U5_Buff_out_reg_2_inst : DF3 port map( D => U5_n25, C => CLK, Q => 
                           Filter_Out(2), QN => U5_n14);
   U5_Buff_out_reg_3_inst : DF3 port map( D => U5_n24, C => CLK, Q => 
                           Filter_Out(3), QN => U5_n15);
   U5_Buff_out_reg_4_inst : DF3 port map( D => U5_n23, C => CLK, Q => 
                           Filter_Out(4), QN => U5_n16);
   U5_Buff_out_reg_5_inst : DF3 port map( D => U5_n22, C => CLK, Q => 
                           Filter_Out(5), QN => U5_n17);
   U5_Buff_out_reg_6_inst : DF3 port map( D => U5_n21, C => CLK, Q => 
                           Filter_Out(6), QN => U5_n18);
   U5_Buff_out_reg_7_inst : DF3 port map( D => U5_n20, C => CLK, Q => 
                           Filter_Out(7), QN => U5_n19);
   U6_U13 : OAI212 port map( A => U6_n33, B => n121, C => n233, Q => U6_n36);
   U6_U6 : OAI212 port map( A => U6_n13, B => U1_n7, C => U6_n29, Q => U6_n42);
   U6_cpt_current_reg_3_inst : DFC3 port map( D => U6_n40, C => CLK, RN => n263
                           , Q => U6_n47, QN => n31);
   U6_cpt_current_reg_2_inst : DFC3 port map( D => U6_n39, C => CLK, RN => n263
                           , Q => n_1139, QN => n19);
   U6_cpt_current_reg_1_inst : DFC3 port map( D => U6_n38, C => CLK, RN => n263
                           , Q => n223, QN => U6_n33);
   U6_cpt_current_reg_4_inst : DFC3 port map( D => U6_n42, C => CLK, RN => n263
                           , Q => U6_n48, QN => n_1140);
   U6_current_state_reg_2_inst : DFC3 port map( D => U6_n41, C => CLK, RN => 
                           n263, Q => n149, QN => U6_n14);
   U6_current_state_reg_1_inst : DFC3 port map( D => U6_n7, C => CLK, RN => 
                           n263, Q => U6_n50, QN => n30);
   U6_cpt_current_reg_0_inst : DFC3 port map( D => U6_n37, C => CLK, RN => n263
                           , Q => U6_n4, QN => n121);
   U6_current_state_reg_0_inst : DFC3 port map( D => U6_n10, C => CLK, RN => 
                           n263, Q => U6_n2, QN => n_1141);
   U7_U10 : OAI212 port map( A => n56, B => n148, C => U7_n12, Q => ADC_Convstb
                           );
   U7_U4 : OAI222 port map( A => U7_n2, B => ack_F2ADC, C => req_ADC2F, D => 
                           U7_n11, Q => U7_n10);
   U7_current_state_reg_1_inst : DFC3 port map( D => U7_n14, C => CLK, RN => 
                           n263, Q => U7_n2, QN => n148);
   U7_current_state_reg_2_inst : DFC3 port map( D => U7_n13, C => CLK, RN => 
                           n263, Q => n56, QN => n_1142);
   U7_current_state_reg_0_inst : DFC3 port map( D => U7_n15, C => CLK, RN => 
                           n263, Q => n150, QN => U7_n9);
   U8_current_state_reg : DF3 port map( D => U8_N5_port, C => CLK, Q => 
                           U8_current_state, QN => DAC_WRb_port);
   U8_pre_req_F2DAC_reg : DF3 port map( D => U8_n1, C => CLK, Q => 
                           U8_pre_req_F2DAC, QN => n_1143);
   U9_U17 : OAI212 port map( A => U9_n1, B => U9_n19, C => U9_n10, Q => U9_n20)
                           ;
   U9_U15 : OAI212 port map( A => U9_n1, B => U9_n18, C => U9_n9, Q => U9_n21);
   U9_U13 : OAI212 port map( A => U9_n1, B => U9_n17, C => U9_n8, Q => U9_n22);
   U9_U11 : OAI212 port map( A => U9_n1, B => U9_n16, C => U9_n7, Q => U9_n23);
   U9_U9 : OAI212 port map( A => U9_n1, B => U9_n15, C => U9_n6, Q => U9_n24);
   U9_U7 : OAI212 port map( A => U9_n1, B => U9_n14, C => U9_n5, Q => U9_n25);
   U9_U5 : OAI212 port map( A => U9_n1, B => U9_n13, C => U9_n4, Q => U9_n26);
   U9_U3 : OAI212 port map( A => U9_n1, B => U9_n12, C => U9_n2, Q => U9_n27);
   U9_reg_reg_0_inst : DF3 port map( D => U9_n27, C => CLK, Q => 
                           Filter_In_mem_0_port, QN => U9_n12);
   U9_reg_reg_1_inst : DF3 port map( D => U9_n26, C => CLK, Q => 
                           Filter_In_mem_1_port, QN => U9_n13);
   U9_reg_reg_2_inst : DF3 port map( D => U9_n25, C => CLK, Q => 
                           Filter_In_mem_2_port, QN => U9_n14);
   U9_reg_reg_3_inst : DF3 port map( D => U9_n24, C => CLK, Q => 
                           Filter_In_mem_3_port, QN => U9_n15);
   U9_reg_reg_4_inst : DF3 port map( D => U9_n23, C => CLK, Q => 
                           Filter_In_mem_4_port, QN => U9_n16);
   U9_reg_reg_5_inst : DF3 port map( D => U9_n22, C => CLK, Q => 
                           Filter_In_mem_5_port, QN => U9_n17);
   U9_reg_reg_6_inst : DF3 port map( D => U9_n21, C => CLK, Q => 
                           Filter_In_mem_6_port, QN => U9_n18);
   U9_reg_reg_7_inst : DF3 port map( D => U9_n20, C => CLK, Q => 
                           Filter_In_mem_7_port, QN => U9_n19);
   U3_mult_19_S3_2_6 : ADD32 port map( A => U3_mult_19_ab_2_6_port, B => 
                           U3_mult_19_CARRYB_1_6_port, CI => 
                           U3_mult_19_ab_1_7_port, CO => 
                           U3_mult_19_CARRYB_2_6_port, S => 
                           U3_mult_19_SUMB_2_6_port);
   U3_mult_19_S2_2_5 : ADD32 port map( A => U3_mult_19_ab_2_5_port, B => 
                           U3_mult_19_CARRYB_1_5_port, CI => 
                           U3_mult_19_SUMB_1_6_port, CO => 
                           U3_mult_19_CARRYB_2_5_port, S => 
                           U3_mult_19_SUMB_2_5_port);
   U3_mult_19_S2_2_4 : ADD32 port map( A => U3_mult_19_ab_2_4_port, B => 
                           U3_mult_19_CARRYB_1_4_port, CI => 
                           U3_mult_19_SUMB_1_5_port, CO => 
                           U3_mult_19_CARRYB_2_4_port, S => 
                           U3_mult_19_SUMB_2_4_port);
   U3_mult_19_S2_2_3 : ADD32 port map( A => U3_mult_19_ab_2_3_port, B => 
                           U3_mult_19_CARRYB_1_3_port, CI => 
                           U3_mult_19_SUMB_1_4_port, CO => 
                           U3_mult_19_CARRYB_2_3_port, S => 
                           U3_mult_19_SUMB_2_3_port);
   U3_mult_19_S2_2_2 : ADD32 port map( A => U3_mult_19_ab_2_2_port, B => 
                           U3_mult_19_CARRYB_1_2_port, CI => 
                           U3_mult_19_SUMB_1_3_port, CO => 
                           U3_mult_19_CARRYB_2_2_port, S => 
                           U3_mult_19_SUMB_2_2_port);
   U3_mult_19_S2_2_1 : ADD32 port map( A => U3_mult_19_ab_2_1_port, B => 
                           U3_mult_19_CARRYB_1_1_port, CI => 
                           U3_mult_19_SUMB_1_2_port, CO => 
                           U3_mult_19_CARRYB_2_1_port, S => 
                           U3_mult_19_SUMB_2_1_port);
   U3_mult_19_S1_2_0 : ADD32 port map( A => U3_mult_19_ab_2_0_port, B => 
                           U3_mult_19_CARRYB_1_0_port, CI => 
                           U3_mult_19_SUMB_1_1_port, CO => 
                           U3_mult_19_CARRYB_2_0_port, S => Mult_out_2_port);
   U3_mult_19_S3_3_6 : ADD32 port map( A => U3_mult_19_ab_3_6_port, B => 
                           U3_mult_19_CARRYB_2_6_port, CI => 
                           U3_mult_19_ab_2_7_port, CO => 
                           U3_mult_19_CARRYB_3_6_port, S => 
                           U3_mult_19_SUMB_3_6_port);
   U3_mult_19_S2_3_5 : ADD32 port map( A => U3_mult_19_ab_3_5_port, B => 
                           U3_mult_19_CARRYB_2_5_port, CI => 
                           U3_mult_19_SUMB_2_6_port, CO => 
                           U3_mult_19_CARRYB_3_5_port, S => 
                           U3_mult_19_SUMB_3_5_port);
   U3_mult_19_S2_3_4 : ADD32 port map( A => U3_mult_19_ab_3_4_port, B => 
                           U3_mult_19_CARRYB_2_4_port, CI => 
                           U3_mult_19_SUMB_2_5_port, CO => 
                           U3_mult_19_CARRYB_3_4_port, S => 
                           U3_mult_19_SUMB_3_4_port);
   U3_mult_19_S2_3_3 : ADD32 port map( A => U3_mult_19_ab_3_3_port, B => 
                           U3_mult_19_CARRYB_2_3_port, CI => 
                           U3_mult_19_SUMB_2_4_port, CO => 
                           U3_mult_19_CARRYB_3_3_port, S => 
                           U3_mult_19_SUMB_3_3_port);
   U3_mult_19_S2_3_2 : ADD32 port map( A => U3_mult_19_ab_3_2_port, B => 
                           U3_mult_19_CARRYB_2_2_port, CI => 
                           U3_mult_19_SUMB_2_3_port, CO => 
                           U3_mult_19_CARRYB_3_2_port, S => 
                           U3_mult_19_SUMB_3_2_port);
   U3_mult_19_S2_3_1 : ADD32 port map( A => U3_mult_19_ab_3_1_port, B => 
                           U3_mult_19_CARRYB_2_1_port, CI => 
                           U3_mult_19_SUMB_2_2_port, CO => 
                           U3_mult_19_CARRYB_3_1_port, S => 
                           U3_mult_19_SUMB_3_1_port);
   U3_mult_19_S1_3_0 : ADD32 port map( A => U3_mult_19_ab_3_0_port, B => 
                           U3_mult_19_CARRYB_2_0_port, CI => 
                           U3_mult_19_SUMB_2_1_port, CO => 
                           U3_mult_19_CARRYB_3_0_port, S => Mult_out_3_port);
   U3_mult_19_S3_4_6 : ADD32 port map( A => U3_mult_19_ab_4_6_port, B => 
                           U3_mult_19_CARRYB_3_6_port, CI => 
                           U3_mult_19_ab_3_7_port, CO => 
                           U3_mult_19_CARRYB_4_6_port, S => 
                           U3_mult_19_SUMB_4_6_port);
   U3_mult_19_S2_4_5 : ADD32 port map( A => U3_mult_19_ab_4_5_port, B => 
                           U3_mult_19_CARRYB_3_5_port, CI => 
                           U3_mult_19_SUMB_3_6_port, CO => 
                           U3_mult_19_CARRYB_4_5_port, S => 
                           U3_mult_19_SUMB_4_5_port);
   U3_mult_19_S2_4_4 : ADD32 port map( A => U3_mult_19_ab_4_4_port, B => 
                           U3_mult_19_CARRYB_3_4_port, CI => 
                           U3_mult_19_SUMB_3_5_port, CO => 
                           U3_mult_19_CARRYB_4_4_port, S => 
                           U3_mult_19_SUMB_4_4_port);
   U3_mult_19_S2_4_3 : ADD32 port map( A => U3_mult_19_ab_4_3_port, B => 
                           U3_mult_19_CARRYB_3_3_port, CI => 
                           U3_mult_19_SUMB_3_4_port, CO => 
                           U3_mult_19_CARRYB_4_3_port, S => 
                           U3_mult_19_SUMB_4_3_port);
   U3_mult_19_S2_4_2 : ADD32 port map( A => U3_mult_19_ab_4_2_port, B => 
                           U3_mult_19_CARRYB_3_2_port, CI => 
                           U3_mult_19_SUMB_3_3_port, CO => 
                           U3_mult_19_CARRYB_4_2_port, S => 
                           U3_mult_19_SUMB_4_2_port);
   U3_mult_19_S2_4_1 : ADD32 port map( A => U3_mult_19_ab_4_1_port, B => 
                           U3_mult_19_CARRYB_3_1_port, CI => 
                           U3_mult_19_SUMB_3_2_port, CO => 
                           U3_mult_19_CARRYB_4_1_port, S => 
                           U3_mult_19_SUMB_4_1_port);
   U3_mult_19_S1_4_0 : ADD32 port map( A => U3_mult_19_ab_4_0_port, B => 
                           U3_mult_19_CARRYB_3_0_port, CI => 
                           U3_mult_19_SUMB_3_1_port, CO => 
                           U3_mult_19_CARRYB_4_0_port, S => Mult_out_4_port);
   U3_mult_19_S3_5_6 : ADD32 port map( A => U3_mult_19_ab_5_6_port, B => 
                           U3_mult_19_CARRYB_4_6_port, CI => 
                           U3_mult_19_ab_4_7_port, CO => 
                           U3_mult_19_CARRYB_5_6_port, S => 
                           U3_mult_19_SUMB_5_6_port);
   U3_mult_19_S2_5_5 : ADD32 port map( A => U3_mult_19_ab_5_5_port, B => 
                           U3_mult_19_CARRYB_4_5_port, CI => 
                           U3_mult_19_SUMB_4_6_port, CO => 
                           U3_mult_19_CARRYB_5_5_port, S => 
                           U3_mult_19_SUMB_5_5_port);
   U3_mult_19_S2_5_4 : ADD32 port map( A => U3_mult_19_ab_5_4_port, B => 
                           U3_mult_19_CARRYB_4_4_port, CI => 
                           U3_mult_19_SUMB_4_5_port, CO => 
                           U3_mult_19_CARRYB_5_4_port, S => 
                           U3_mult_19_SUMB_5_4_port);
   U3_mult_19_S2_5_3 : ADD32 port map( A => U3_mult_19_ab_5_3_port, B => 
                           U3_mult_19_CARRYB_4_3_port, CI => 
                           U3_mult_19_SUMB_4_4_port, CO => 
                           U3_mult_19_CARRYB_5_3_port, S => 
                           U3_mult_19_SUMB_5_3_port);
   U3_mult_19_S2_5_2 : ADD32 port map( A => U3_mult_19_ab_5_2_port, B => 
                           U3_mult_19_CARRYB_4_2_port, CI => 
                           U3_mult_19_SUMB_4_3_port, CO => 
                           U3_mult_19_CARRYB_5_2_port, S => 
                           U3_mult_19_SUMB_5_2_port);
   U3_mult_19_S2_5_1 : ADD32 port map( A => U3_mult_19_ab_5_1_port, B => 
                           U3_mult_19_CARRYB_4_1_port, CI => 
                           U3_mult_19_SUMB_4_2_port, CO => 
                           U3_mult_19_CARRYB_5_1_port, S => 
                           U3_mult_19_SUMB_5_1_port);
   U3_mult_19_S1_5_0 : ADD32 port map( A => U3_mult_19_ab_5_0_port, B => 
                           U3_mult_19_CARRYB_4_0_port, CI => 
                           U3_mult_19_SUMB_4_1_port, CO => 
                           U3_mult_19_CARRYB_5_0_port, S => Mult_out_5_port);
   U3_mult_19_S3_6_6 : ADD32 port map( A => U3_mult_19_ab_6_6_port, B => 
                           U3_mult_19_CARRYB_5_6_port, CI => 
                           U3_mult_19_ab_5_7_port, CO => 
                           U3_mult_19_CARRYB_6_6_port, S => 
                           U3_mult_19_SUMB_6_6_port);
   U3_mult_19_S2_6_5 : ADD32 port map( A => U3_mult_19_ab_6_5_port, B => 
                           U3_mult_19_CARRYB_5_5_port, CI => 
                           U3_mult_19_SUMB_5_6_port, CO => 
                           U3_mult_19_CARRYB_6_5_port, S => 
                           U3_mult_19_SUMB_6_5_port);
   U3_mult_19_S2_6_4 : ADD32 port map( A => U3_mult_19_ab_6_4_port, B => 
                           U3_mult_19_CARRYB_5_4_port, CI => 
                           U3_mult_19_SUMB_5_5_port, CO => 
                           U3_mult_19_CARRYB_6_4_port, S => 
                           U3_mult_19_SUMB_6_4_port);
   U3_mult_19_S2_6_3 : ADD32 port map( A => U3_mult_19_ab_6_3_port, B => 
                           U3_mult_19_CARRYB_5_3_port, CI => 
                           U3_mult_19_SUMB_5_4_port, CO => 
                           U3_mult_19_CARRYB_6_3_port, S => 
                           U3_mult_19_SUMB_6_3_port);
   U3_mult_19_S2_6_2 : ADD32 port map( A => U3_mult_19_ab_6_2_port, B => 
                           U3_mult_19_CARRYB_5_2_port, CI => 
                           U3_mult_19_SUMB_5_3_port, CO => 
                           U3_mult_19_CARRYB_6_2_port, S => 
                           U3_mult_19_SUMB_6_2_port);
   U3_mult_19_S2_6_1 : ADD32 port map( A => U3_mult_19_ab_6_1_port, B => 
                           U3_mult_19_CARRYB_5_1_port, CI => 
                           U3_mult_19_SUMB_5_2_port, CO => 
                           U3_mult_19_CARRYB_6_1_port, S => 
                           U3_mult_19_SUMB_6_1_port);
   U3_mult_19_S1_6_0 : ADD32 port map( A => U3_mult_19_ab_6_0_port, B => 
                           U3_mult_19_CARRYB_5_0_port, CI => 
                           U3_mult_19_SUMB_5_1_port, CO => 
                           U3_mult_19_CARRYB_6_0_port, S => Mult_out_6_port);
   U3_mult_19_S5_6 : ADD32 port map( A => U3_mult_19_ab_7_6_port, B => 
                           U3_mult_19_CARRYB_6_6_port, CI => 
                           U3_mult_19_ab_6_7_port, CO => 
                           U3_mult_19_CARRYB_7_6_port, S => 
                           U3_mult_19_SUMB_7_6_port);
   U3_mult_19_S4_5 : ADD32 port map( A => U3_mult_19_ab_7_5_port, B => 
                           U3_mult_19_CARRYB_6_5_port, CI => 
                           U3_mult_19_SUMB_6_6_port, CO => 
                           U3_mult_19_CARRYB_7_5_port, S => 
                           U3_mult_19_SUMB_7_5_port);
   U3_mult_19_S4_4 : ADD32 port map( A => U3_mult_19_ab_7_4_port, B => 
                           U3_mult_19_CARRYB_6_4_port, CI => 
                           U3_mult_19_SUMB_6_5_port, CO => 
                           U3_mult_19_CARRYB_7_4_port, S => 
                           U3_mult_19_SUMB_7_4_port);
   U3_mult_19_S4_3 : ADD32 port map( A => U3_mult_19_ab_7_3_port, B => 
                           U3_mult_19_CARRYB_6_3_port, CI => 
                           U3_mult_19_SUMB_6_4_port, CO => 
                           U3_mult_19_CARRYB_7_3_port, S => 
                           U3_mult_19_SUMB_7_3_port);
   U3_mult_19_S4_2 : ADD32 port map( A => U3_mult_19_ab_7_2_port, B => 
                           U3_mult_19_CARRYB_6_2_port, CI => 
                           U3_mult_19_SUMB_6_3_port, CO => 
                           U3_mult_19_CARRYB_7_2_port, S => 
                           U3_mult_19_SUMB_7_2_port);
   U3_mult_19_S4_1 : ADD32 port map( A => U3_mult_19_ab_7_1_port, B => 
                           U3_mult_19_CARRYB_6_1_port, CI => 
                           U3_mult_19_SUMB_6_2_port, CO => 
                           U3_mult_19_CARRYB_7_1_port, S => 
                           U3_mult_19_SUMB_7_1_port);
   U3_mult_19_S4_0 : ADD32 port map( A => U3_mult_19_ab_7_0_port, B => 
                           U3_mult_19_CARRYB_6_0_port, CI => 
                           U3_mult_19_SUMB_6_1_port, CO => 
                           U3_mult_19_CARRYB_7_0_port, S => Mult_out_7_port);
   U4_add_27_aco_U1_1 : ADD32 port map( A => U4_N49, B => Mult_out_1_port, CI 
                           => U4_add_27_aco_carry_1_port, CO => 
                           U4_add_27_aco_carry_2_port, S => U4_N7);
   U4_add_27_aco_U1_2 : ADD32 port map( A => U4_N50, B => Mult_out_2_port, CI 
                           => U4_add_27_aco_carry_2_port, CO => 
                           U4_add_27_aco_carry_3_port, S => U4_N8);
   U4_add_27_aco_U1_3 : ADD32 port map( A => U4_N51, B => Mult_out_3_port, CI 
                           => U4_add_27_aco_carry_3_port, CO => 
                           U4_add_27_aco_carry_4_port, S => U4_N9);
   U4_add_27_aco_U1_4 : ADD32 port map( A => U4_N52, B => Mult_out_4_port, CI 
                           => U4_add_27_aco_carry_4_port, CO => 
                           U4_add_27_aco_carry_5_port, S => U4_N10);
   U4_add_27_aco_U1_5 : ADD32 port map( A => U4_N53, B => Mult_out_5_port, CI 
                           => U4_add_27_aco_carry_5_port, CO => 
                           U4_add_27_aco_carry_6_port, S => U4_N11);
   U4_add_27_aco_U1_6 : ADD32 port map( A => U4_N54, B => Mult_out_6_port, CI 
                           => U4_add_27_aco_carry_6_port, CO => 
                           U4_add_27_aco_carry_7_port, S => U4_N12);
   U4_add_27_aco_U1_7 : ADD32 port map( A => U4_N55, B => Mult_out_7_port, CI 
                           => U4_add_27_aco_carry_7_port, CO => 
                           U4_add_27_aco_carry_8_port, S => U4_N13);
   U4_add_27_aco_U1_8 : ADD32 port map( A => U4_N56, B => Mult_out_8_port, CI 
                           => U4_add_27_aco_carry_8_port, CO => 
                           U4_add_27_aco_carry_9_port, S => U4_N14);
   U4_add_27_aco_U1_9 : ADD32 port map( A => U4_N57, B => Mult_out_9_port, CI 
                           => U4_add_27_aco_carry_9_port, CO => 
                           U4_add_27_aco_carry_10_port, S => U4_N15);
   U4_add_27_aco_U1_10 : ADD32 port map( A => U4_N58, B => Mult_out_10_port, CI
                           => U4_add_27_aco_carry_10_port, CO => 
                           U4_add_27_aco_carry_11_port, S => U4_N16);
   U4_add_27_aco_U1_11 : ADD32 port map( A => U4_N59, B => Mult_out_11_port, CI
                           => U4_add_27_aco_carry_11_port, CO => 
                           U4_add_27_aco_carry_12_port, S => U4_N17);
   U4_add_27_aco_U1_12 : ADD32 port map( A => U4_N60, B => Mult_out_12_port, CI
                           => U4_add_27_aco_carry_12_port, CO => 
                           U4_add_27_aco_carry_13_port, S => U4_N18);
   U4_add_27_aco_U1_13 : ADD32 port map( A => U4_N61, B => Mult_out_13_port, CI
                           => U4_add_27_aco_carry_13_port, CO => 
                           U4_add_27_aco_carry_14_port, S => U4_N19);
   U4_add_27_aco_U1_14 : ADD32 port map( A => U4_N62, B => Mult_out_14_port, CI
                           => U4_add_27_aco_carry_14_port, CO => 
                           U4_add_27_aco_carry_15_port, S => U4_N20);
   U4_add_27_aco_U1_15 : ADD32 port map( A => U4_N63, B => Mult_out_15_port, CI
                           => U4_add_27_aco_carry_15_port, CO => 
                           U4_add_27_aco_carry_16_port, S => U4_N21);
   U3_mult_19_FS_1_U37 : OAI212 port map( A => U3_mult_19_FS_1_n12, B => 
                           U3_mult_19_FS_1_n31, C => U3_mult_19_FS_1_n13, Q => 
                           U3_mult_19_FS_1_n9);
   U3_mult_19_FS_1_U28 : XOR31 port map( A => U3_mult_19_A2_11_port, B => 
                           U3_mult_19_A1_11_port, C => U3_mult_19_FS_1_n28, Q 
                           => Mult_out_13_port);
   U3_mult_19_FS_1_U27 : OAI212 port map( A => U3_mult_19_FS_1_n13, B => 
                           U3_mult_19_FS_1_n22, C => U3_mult_19_FS_1_n11, Q => 
                           U3_mult_19_FS_1_n27);
   U3_mult_19_FS_1_U26 : OAI212 port map( A => U3_mult_19_FS_1_n23, B => 
                           U3_mult_19_FS_1_n37, C => U3_mult_19_FS_1_n26, Q => 
                           U3_mult_19_FS_1_n20);
   U3_mult_19_FS_1_U25 : OAI212 port map( A => U3_mult_19_A1_11_port, B => 
                           U3_mult_19_FS_1_n20, C => U3_mult_19_A2_11_port, Q 
                           => U3_mult_19_FS_1_n25);
   U3_mult_19_FS_1_U21 : XOR31 port map( A => U3_mult_19_A2_12_port, B => 
                           U3_mult_19_A1_12_port, C => U3_mult_19_FS_1_n33, Q 
                           => Mult_out_14_port);
   U3_mult_19_FS_1_U20 : OAI212 port map( A => U3_mult_19_A1_12_port, B => 
                           U3_mult_19_FS_1_n33, C => U3_mult_19_A2_12_port, Q 
                           => U3_mult_19_FS_1_n18);
   U3_mult_19_FS_1_U15 : OAI212 port map( A => U3_mult_19_FS_1_n12, B => 
                           U3_mult_19_FS_1_n13, C => U3_mult_19_FS_1_n14, Q => 
                           Mult_out_10_port);
   U12 : NOR22 port map( A => U6_n44, B => U6_n33, Q => n229);
   U13 : NAND22 port map( A => U3_mult_19_ab_0_2_port, B => 
                           U3_mult_19_ab_1_1_port, Q => n3);
   U14 : INV3 port map( A => n3, Q => U3_mult_19_CARRYB_1_1_port);
   U15 : MUX22 port map( A => U2_n523, B => U2_n522, S => U6_n29, Q => 
                           U3_mult_19_n64);
   U16 : NAND22 port map( A => U3_mult_19_CARRYB_7_3_port, B => 
                           U3_mult_19_SUMB_7_4_port, Q => n4);
   U17 : INV3 port map( A => n4, Q => U3_mult_19_A2_10_port);
   U18 : NOR30 port map( A => n149, B => U6_n2, C => n30, Q => Buff_OE);
   U19 : MUX22 port map( A => U2_n613, B => U2_n612, S => U6_n29, Q => 
                           U3_mult_19_n65);
   U20 : NAND22 port map( A => U3_mult_19_CARRYB_7_4_port, B => 
                           U3_mult_19_SUMB_7_5_port, Q => n5);
   U21 : INV3 port map( A => n5, Q => U3_mult_19_A2_11_port);
   U22 : NOR20 port map( A => U6_n16, B => U6_n2, Q => Delay_Line_sample_shift)
                           ;
   U23 : XNR21 port map( A => n11, B => U3_mult_19_A1_7_port, Q => 
                           Mult_out_9_port);
   U24 : NAND22 port map( A => U3_mult_19_ab_0_7_port, B => 
                           U3_mult_19_ab_1_6_port, Q => n6);
   U25 : INV3 port map( A => n6, Q => U3_mult_19_CARRYB_1_6_port);
   U26 : XNR31 port map( A => U3_mult_19_FS_1_n29, B => U3_mult_19_A2_10_port, 
                           C => U3_mult_19_A1_10_port, Q => Mult_out_12_port);
   U27 : NAND22 port map( A => U3_mult_19_CARRYB_7_1_port, B => 
                           U3_mult_19_SUMB_7_2_port, Q => n7);
   U28 : INV3 port map( A => n7, Q => U3_mult_19_A2_8_port);
   U29 : MUX22 port map( A => U2_n701, B => U2_n700, S => U6_n29, Q => 
                           U3_mult_19_n83);
   U30 : AOI211 port map( A => U6_n2, B => ack_F2ADC, C => n8, Q => U4_N61);
   U31 : MUX22 port map( A => U2_n351, B => U2_n350, S => U6_n29, Q => 
                           U3_mult_19_n62);
   U32 : NAND22 port map( A => U3_mult_19_ab_0_1_port, B => 
                           U3_mult_19_ab_1_0_port, Q => n9);
   U33 : INV3 port map( A => n9, Q => U3_mult_19_CARRYB_1_0_port);
   U34 : XOR21 port map( A => U3_mult_19_FS_1_n17, B => n13, Q => 
                           Mult_out_15_port);
   U35 : NAND22 port map( A => U3_mult_19_ab_0_6_port, B => 
                           U3_mult_19_ab_1_5_port, Q => n10);
   U36 : INV3 port map( A => n10, Q => U3_mult_19_CARRYB_1_5_port);
   U37 : AOI311 port map( A => n56, B => U7_n9, C => n148, D => RESET, Q => 
                           U9_n11);
   U38 : NAND22 port map( A => U3_mult_19_CARRYB_7_0_port, B => 
                           U3_mult_19_SUMB_7_1_port, Q => n11);
   U39 : INV3 port map( A => n11, Q => U3_mult_19_A2_7_port);
   U40 : OAI212 port map( A => U3_mult_19_A2_9_port, B => U3_mult_19_A1_9_port,
                           C => U3_mult_19_FS_1_n11, Q => U3_mult_19_FS_1_n10);
   U41 : NAND22 port map( A => U3_mult_19_CARRYB_7_5_port, B => 
                           U3_mult_19_SUMB_7_6_port, Q => n12);
   U42 : INV3 port map( A => n12, Q => U3_mult_19_A2_12_port);
   U43 : NOR31 port map( A => U4_add_27_aco_n18, B => 
                           U4_mult_add_27_aco_PROD_not_16_port, C => 
                           U4_mult_add_27_aco_PROD_not_17_port, Q => 
                           U4_add_27_aco_carry_18_port);
   U44 : IMUX21 port map( A => U1_n51, B => U1_n18, S => Rom_Address_2_port, Q 
                           => U1_n48);
   U45 : IMAJ31 port map( A => U3_mult_19_FS_1_n9, B => U3_mult_19_A2_9_port, C
                           => U3_mult_19_A1_9_port, Q => U3_mult_19_FS_1_n29);
   U46 : NAND22 port map( A => U3_mult_19_CARRYB_7_6_port, B => 
                           U3_mult_19_ab_7_7_port, Q => n13);
   U47 : AOI211 port map( A => U6_n31, B => req_ADC2F, C => 
                           Delay_Line_sample_shift, Q => n14);
   U48 : INV3 port map( A => n14, Q => U6_n41);
   U49 : XOR21 port map( A => U4_mult_add_27_aco_PROD_not_0_port, B => 
                           Mult_out_0_port, Q => n228);
   U50 : NOR21 port map( A => RESET, B => n228, Q => U4_N27);
   U51 : NOR21 port map( A => RESET, B => n225, Q => U4_N43);
   U52 : NOR21 port map( A => RESET, B => n226, Q => U4_N44);
   U53 : NOR21 port map( A => RESET, B => n227, Q => U4_N45);
   U54 : NOR21 port map( A => n232, B => n231, Q => U2_n716);
   U55 : NAND22 port map( A => U2_n716, B => U2_n717, Q => U2_n357);
   U56 : NAND22 port map( A => U2_n716, B => U2_n720, Q => U2_n358);
   U57 : CLKIN3 port map( A => n230, Q => U1_n12);
   U58 : INV3 port map( A => n229, Q => U2_n280);
   U59 : INV3 port map( A => U2_n723, Q => U2_n269);
   U60 : BUF2 port map( A => Rom_Address_0_port, Q => n230);
   U61 : XOR21 port map( A => U4_mult_add_27_aco_PROD_not_19_port, B => 
                           U4_add_27_aco_carry_19_port, Q => n224);
   U62 : NAND22 port map( A => U3_mult_19_A2_8_port, B => U3_mult_19_A1_8_port,
                           Q => U3_mult_19_FS_1_n13);
   U63 : NAND20 port map( A => U2_n718, B => U2_n724, Q => U2_n726);
   U64 : INV1 port map( A => U3_mult_19_ab_1_2_port, Q => U3_mult_19_n70);
   U65 : INV2 port map( A => U3_mult_19_ab_0_4_port, Q => U3_mult_19_n79);
   U66 : NAND22 port map( A => U2_n716, B => U2_n719, Q => U2_n359);
   U67 : INV3 port map( A => U2_n734, Q => U2_n276);
   U68 : CLKIN1 port map( A => n231, Q => U2_n278);
   U69 : INV3 port map( A => U4_add_27_aco_carry_16_port, Q => 
                           U4_add_27_aco_n18);
   U70 : OAI222 port map( A => n15, B => U2_n358, C => n32, D => U2_n359, Q => 
                           U2_n682);
   U71 : INV3 port map( A => Delay_Line_out_1_port, Q => U3_mult_19_n75);
   U72 : AOI221 port map( A => U2_n272, B => U2_x_12_1_port, C => U2_n273, D =>
                           U2_x_13_1_port, Q => U2_n697);
   U73 : AOI221 port map( A => U2_n274, B => U2_x_10_1_port, C => U2_n275, D =>
                           U2_x_11_1_port, Q => U2_n698);
   U74 : AOI221 port map( A => U2_n276, B => U2_x_8_1_port, C => U2_n277, D => 
                           U2_x_9_1_port, Q => U2_n699);
   U75 : NOR20 port map( A => n121, B => U6_n44, Q => Rom_Address_0_port);
   U76 : OAI211 port map( A => U3_mult_19_FS_1_n23, B => U3_mult_19_FS_1_n29, C
                           => U3_mult_19_FS_1_n26, Q => U3_mult_19_FS_1_n28);
   U77 : NOR20 port map( A => U3_mult_19_A1_8_port, B => U3_mult_19_A2_8_port, 
                           Q => U3_mult_19_FS_1_n31);
   U78 : NOR20 port map( A => U3_mult_19_A1_8_port, B => U3_mult_19_FS_1_n39, Q
                           => U3_mult_19_FS_1_n16);
   U79 : INV1 port map( A => U3_mult_19_FS_1_n12, Q => U3_mult_19_FS_1_n39);
   U80 : OAI220 port map( A => U3_mult_19_A1_11_port, B => 
                           U3_mult_19_A2_11_port, C => U3_mult_19_A1_8_port, D 
                           => U3_mult_19_A2_8_port, Q => U3_mult_19_FS_1_n24);
   U81 : NAND20 port map( A => U2_n717, B => U2_n724, Q => U2_n727);
   U82 : CLKIN3 port map( A => U2_n741, Q => U2_n270);
   U83 : NAND21 port map( A => U2_n738, B => U2_n717, Q => U2_n741);
   U84 : CLKIN3 port map( A => U2_n725, Q => U2_n268);
   U85 : NAND20 port map( A => U2_n724, B => U2_n719, Q => U2_n725);
   U86 : NAND20 port map( A => U2_n720, B => U2_n724, Q => U2_n723);
   U87 : CLKIN3 port map( A => U2_n737, Q => U2_n273);
   U88 : NAND21 port map( A => U2_n738, B => U2_n720, Q => U2_n737);
   U89 : NOR20 port map( A => U3_mult_19_n88, B => U3_mult_19_n75, Q => 
                           U3_mult_19_ab_1_3_port);
   U90 : NOR20 port map( A => U3_mult_19_n90, B => U3_mult_19_n75, Q => 
                           U3_mult_19_ab_1_1_port);
   U91 : NOR20 port map( A => U3_mult_19_n91, B => U3_mult_19_n75, Q => 
                           U3_mult_19_ab_1_0_port);
   U92 : NOR20 port map( A => U3_mult_19_n89, B => U3_mult_19_n75, Q => 
                           U3_mult_19_ab_1_2_port);
   U93 : NOR20 port map( A => U3_mult_19_n89, B => U3_mult_19_n83, Q => 
                           U3_mult_19_ab_0_2_port);
   U94 : NOR20 port map( A => U3_mult_19_n90, B => U3_mult_19_n83, Q => 
                           U3_mult_19_ab_0_1_port);
   U95 : NOR20 port map( A => U3_mult_19_n88, B => U3_mult_19_n83, Q => 
                           U3_mult_19_ab_0_3_port);
   U96 : NOR20 port map( A => U3_mult_19_n87, B => U3_mult_19_n83, Q => 
                           U3_mult_19_ab_0_4_port);
   U97 : NOR20 port map( A => U3_mult_19_n84, B => U3_mult_19_n75, Q => 
                           U3_mult_19_ab_1_7_port);
   U98 : INV2 port map( A => n231, Q => U1_n7);
   U99 : NAND21 port map( A => Rom_Address_4_port, B => n231, Q => U1_n20);
   U100 : NOR20 port map( A => U1_n40, B => n231, Q => U1_n28);
   U101 : NAND30 port map( A => Rom_Address_4_port, B => U2_n280, C => n230, Q 
                           => U1_n26);
   U102 : AOI220 port map( A => U1_n23, B => U1_n7, C => U1_n24, D => n230, Q 
                           => U1_n22);
   U103 : OAI210 port map( A => n231, B => Rom_Address_4_port, C => U1_n20, Q 
                           => U1_n37);
   U104 : NAND20 port map( A => n230, B => n233, Q => U1_n30);
   U105 : OAI210 port map( A => n230, B => U1_n25, C => U1_n26, Q => U1_n23);
   U106 : NOR20 port map( A => U3_mult_19_n91, B => U3_mult_19_n83, Q => 
                           Mult_out_0_port);
   U107 : AOI210 port map( A => n230, B => U2_n280, C => U1_n20, Q => U1_n43);
   U108 : OAI310 port map( A => U2_n280, B => n231, C => U1_n2, D => U1_n26, Q 
                           => U1_n50);
   U109 : NAND20 port map( A => U2_n733, B => U2_n719, Q => U2_n734);
   U110 : OAI221 port map( A => n125, B => U2_n358, C => n35, D => U2_n359, Q 
                           => U2_n714);
   U111 : OAI221 port map( A => n127, B => U2_n358, C => n37, D => U2_n359, Q 
                           => U2_n704);
   U112 : OAI220 port map( A => n130, B => U2_n358, C => n40, D => U2_n359, Q 
                           => U2_n660);
   U113 : OAI220 port map( A => n128, B => U2_n358, C => n38, D => U2_n359, Q 
                           => U2_n670);
   U114 : OAI221 port map( A => n126, B => U2_n356, C => n36, D => n235, Q => 
                           U2_n715);
   U115 : OAI221 port map( A => n21, B => U2_n356, C => n16, D => n235, Q => 
                           U2_n705);
   U116 : OAI221 port map( A => n20, B => U2_n356, C => n124, D => n235, Q => 
                           U2_n683);
   U117 : OAI220 port map( A => n22, B => U2_n356, C => n41, D => n235, Q => 
                           U2_n661);
   U118 : OAI220 port map( A => n129, B => U2_n356, C => n39, D => n235, Q => 
                           U2_n671);
   U119 : XNR20 port map( A => U4_N65, B => U4_add_27_aco_carry_17_port, Q => 
                           n226);
   U120 : XNR20 port map( A => U4_N66, B => U4_add_27_aco_carry_18_port, Q => 
                           n227);
   U121 : OAI211 port map( A => n229, B => U1_n12, C => U1_n29, Q => U1_n32);
   U122 : NAND21 port map( A => n229, B => U1_n12, Q => U1_n29);
   U123 : NAND20 port map( A => n229, B => n230, Q => U1_n40);
   U124 : OAI220 port map( A => n133, B => U2_n358, C => n44, D => U2_n359, Q 
                           => U2_n638);
   U125 : OAI220 port map( A => n131, B => U2_n358, C => n42, D => U2_n359, Q 
                           => U2_n648);
   U126 : OAI220 port map( A => n23, B => U2_n356, C => n45, D => n235, Q => 
                           U2_n639);
   U127 : OAI220 port map( A => n132, B => U2_n356, C => n43, D => n235, Q => 
                           U2_n649);
   U128 : XNR20 port map( A => U4_N64, B => U4_add_27_aco_carry_16_port, Q => 
                           n225);
   U129 : OAI210 port map( A => n229, B => U1_n7, C => U1_n29, Q => U1_n51);
   U130 : AOI220 port map( A => U2_n270, B => U2_x_14_1_port, C => U2_n271, D 
                           => U2_x_15_1_port, Q => U2_n696);
   U131 : AOI220 port map( A => U2_n274, B => U2_x_10_0_port, C => U2_n275, D 
                           => U2_x_11_0_port, Q => U2_n730);
   U132 : AOI220 port map( A => U2_n276, B => U2_x_8_0_port, C => U2_n277, D =>
                           U2_x_9_0_port, Q => U2_n731);
   U133 : AOI220 port map( A => U2_n270, B => U2_x_14_0_port, C => U2_n271, D 
                           => U2_x_15_0_port, Q => U2_n728);
   U134 : AOI220 port map( A => U2_n274, B => U2_x_26_2_port, C => U2_n275, D 
                           => U2_x_27_2_port, Q => U2_n666);
   U135 : AOI220 port map( A => U2_n276, B => U2_x_24_2_port, C => U2_n277, D 
                           => U2_x_25_2_port, Q => U2_n667);
   U136 : AOI220 port map( A => U2_n270, B => U2_x_30_2_port, C => U2_n271, D 
                           => U2_x_31_2_port, Q => U2_n664);
   U137 : AOI220 port map( A => U2_n276, B => U2_x_8_2_port, C => U2_n277, D =>
                           U2_x_9_2_port, Q => U2_n677);
   U138 : AOI220 port map( A => U2_n274, B => U2_x_10_2_port, C => U2_n275, D 
                           => U2_x_11_2_port, Q => U2_n676);
   U139 : AOI220 port map( A => U2_n270, B => U2_x_14_2_port, C => U2_n271, D 
                           => U2_x_15_2_port, Q => U2_n674);
   U140 : AOI220 port map( A => U2_n274, B => U2_x_26_3_port, C => U2_n275, D 
                           => U2_x_27_3_port, Q => U2_n644);
   U141 : AOI220 port map( A => U2_n276, B => U2_x_24_3_port, C => U2_n277, D 
                           => U2_x_25_3_port, Q => U2_n645);
   U142 : AOI220 port map( A => U2_n270, B => U2_x_30_3_port, C => U2_n271, D 
                           => U2_x_31_3_port, Q => U2_n642);
   U143 : AOI220 port map( A => U2_n274, B => U2_x_10_3_port, C => U2_n275, D 
                           => U2_x_11_3_port, Q => U2_n654);
   U144 : AOI220 port map( A => U2_n276, B => U2_x_8_3_port, C => U2_n277, D =>
                           U2_x_9_3_port, Q => U2_n655);
   U145 : AOI220 port map( A => U2_n270, B => U2_x_14_3_port, C => U2_n271, D 
                           => U2_x_15_3_port, Q => U2_n652);
   U146 : AOI220 port map( A => U2_n272, B => U2_x_12_0_port, C => U2_n273, D 
                           => U2_x_13_0_port, Q => U2_n729);
   U147 : AOI220 port map( A => U2_n272, B => U2_x_28_2_port, C => U2_n273, D 
                           => U2_x_29_2_port, Q => U2_n665);
   U148 : AOI220 port map( A => U2_n272, B => U2_x_12_2_port, C => U2_n273, D 
                           => U2_x_13_2_port, Q => U2_n675);
   U149 : AOI220 port map( A => U2_n272, B => U2_x_28_3_port, C => U2_n273, D 
                           => U2_x_29_3_port, Q => U2_n643);
   U150 : AOI220 port map( A => U2_n272, B => U2_x_12_3_port, C => U2_n273, D 
                           => U2_x_13_3_port, Q => U2_n653);
   U151 : XOR20 port map( A => U3_mult_19_SUMB_7_1_port, B => 
                           U3_mult_19_CARRYB_7_0_port, Q => Mult_out_8_port);
   U152 : AOI220 port map( A => U2_n268, B => U2_x_0_1_port, C => U2_n269, D =>
                           U2_x_1_1_port, Q => U2_n695);
   U153 : AOI220 port map( A => U2_n268, B => U2_x_0_0_port, C => U2_n269, D =>
                           U2_x_1_0_port, Q => U2_n722);
   U154 : AOI220 port map( A => U2_n266, B => U2_x_18_2_port, C => U2_n267, D 
                           => U2_x_19_2_port, Q => U2_n662);
   U155 : AOI220 port map( A => U2_n268, B => U2_x_16_2_port, C => U2_n269, D 
                           => U2_x_17_2_port, Q => U2_n663);
   U156 : AOI220 port map( A => U2_n268, B => U2_x_0_2_port, C => U2_n269, D =>
                           U2_x_1_2_port, Q => U2_n673);
   U157 : AOI220 port map( A => U2_n266, B => U2_x_2_2_port, C => U2_n267, D =>
                           U2_x_3_2_port, Q => U2_n672);
   U158 : AOI220 port map( A => U2_n266, B => U2_x_18_3_port, C => U2_n267, D 
                           => U2_x_19_3_port, Q => U2_n640);
   U159 : AOI220 port map( A => U2_n268, B => U2_x_16_3_port, C => U2_n269, D 
                           => U2_x_17_3_port, Q => U2_n641);
   U160 : AOI220 port map( A => U2_n274, B => U2_x_26_4_port, C => U2_n275, D 
                           => U2_x_27_4_port, Q => U2_n622);
   U161 : AOI220 port map( A => U2_n276, B => U2_x_24_4_port, C => U2_n277, D 
                           => U2_x_25_4_port, Q => U2_n623);
   U162 : AOI220 port map( A => U2_n270, B => U2_x_30_4_port, C => U2_n271, D 
                           => U2_x_31_4_port, Q => U2_n620);
   U163 : AOI220 port map( A => U2_n274, B => U2_x_10_4_port, C => U2_n275, D 
                           => U2_x_11_4_port, Q => U2_n632);
   U164 : AOI220 port map( A => U2_n276, B => U2_x_8_4_port, C => U2_n277, D =>
                           U2_x_9_4_port, Q => U2_n633);
   U165 : AOI220 port map( A => U2_n270, B => U2_x_14_4_port, C => U2_n271, D 
                           => U2_x_15_4_port, Q => U2_n630);
   U166 : AOI220 port map( A => U2_n274, B => U2_x_26_5_port, C => U2_n275, D 
                           => U2_x_27_5_port, Q => U2_n600);
   U167 : AOI220 port map( A => U2_n276, B => U2_x_24_5_port, C => U2_n277, D 
                           => U2_x_25_5_port, Q => U2_n601);
   U168 : AOI220 port map( A => U2_n270, B => U2_x_30_5_port, C => U2_n271, D 
                           => U2_x_31_5_port, Q => U2_n598);
   U169 : AOI220 port map( A => U2_n274, B => U2_x_10_5_port, C => U2_n275, D 
                           => U2_x_11_5_port, Q => U2_n610);
   U170 : AOI220 port map( A => U2_n276, B => U2_x_8_5_port, C => U2_n277, D =>
                           U2_x_9_5_port, Q => U2_n611);
   U171 : AOI220 port map( A => U2_n270, B => U2_x_14_5_port, C => U2_n271, D 
                           => U2_x_15_5_port, Q => U2_n608);
   U172 : AOI220 port map( A => U2_n266, B => U2_x_18_5_port, C => U2_n267, D 
                           => U2_x_19_5_port, Q => U2_n596);
   U173 : AOI220 port map( A => U2_n268, B => U2_x_16_5_port, C => U2_n269, D 
                           => U2_x_17_5_port, Q => U2_n597);
   U174 : AOI220 port map( A => U2_n272, B => U2_x_28_4_port, C => U2_n273, D 
                           => U2_x_29_4_port, Q => U2_n621);
   U175 : AOI220 port map( A => U2_n272, B => U2_x_12_4_port, C => U2_n273, D 
                           => U2_x_13_4_port, Q => U2_n631);
   U176 : AOI220 port map( A => U2_n272, B => U2_x_28_5_port, C => U2_n273, D 
                           => U2_x_29_5_port, Q => U2_n599);
   U177 : AOI220 port map( A => U2_n272, B => U2_x_12_5_port, C => U2_n273, D 
                           => U2_x_13_5_port, Q => U2_n609);
   U178 : AOI220 port map( A => U2_n266, B => U2_x_2_3_port, C => U2_n267, D =>
                           U2_x_3_3_port, Q => U2_n650);
   U179 : AOI220 port map( A => U2_n268, B => U2_x_0_3_port, C => U2_n269, D =>
                           U2_x_1_3_port, Q => U2_n651);
   U180 : AOI220 port map( A => U2_n266, B => U2_x_18_4_port, C => U2_n267, D 
                           => U2_x_19_4_port, Q => U2_n618);
   U181 : AOI220 port map( A => U2_n268, B => U2_x_16_4_port, C => U2_n269, D 
                           => U2_x_17_4_port, Q => U2_n619);
   U182 : AOI220 port map( A => U2_n266, B => U2_x_2_4_port, C => U2_n267, D =>
                           U2_x_3_4_port, Q => U2_n628);
   U183 : AOI220 port map( A => U2_n268, B => U2_x_0_4_port, C => U2_n269, D =>
                           U2_x_1_4_port, Q => U2_n629);
   U184 : AOI220 port map( A => U2_n266, B => U2_x_2_5_port, C => U2_n267, D =>
                           U2_x_3_5_port, Q => U2_n606);
   U185 : AOI220 port map( A => U2_n268, B => U2_x_0_5_port, C => U2_n269, D =>
                           U2_x_1_5_port, Q => U2_n607);
   U186 : AOI220 port map( A => U2_n266, B => U2_x_18_6_port, C => U2_n267, D 
                           => U2_x_19_6_port, Q => U2_n382);
   U187 : AOI220 port map( A => U2_n268, B => U2_x_16_6_port, C => U2_n269, D 
                           => U2_x_17_6_port, Q => U2_n383);
   U188 : AOI220 port map( A => U2_n266, B => U2_x_2_6_port, C => U2_n267, D =>
                           U2_x_3_6_port, Q => U2_n516);
   U189 : AOI220 port map( A => U2_n268, B => U2_x_0_6_port, C => U2_n269, D =>
                           U2_x_1_6_port, Q => U2_n517);
   U190 : AOI220 port map( A => U2_n274, B => U2_x_26_6_port, C => U2_n275, D 
                           => U2_x_27_6_port, Q => U2_n386);
   U191 : AOI220 port map( A => U2_n276, B => U2_x_24_6_port, C => U2_n277, D 
                           => U2_x_25_6_port, Q => U2_n387);
   U192 : AOI220 port map( A => U2_n270, B => U2_x_30_6_port, C => U2_n271, D 
                           => U2_x_31_6_port, Q => U2_n384);
   U193 : AOI220 port map( A => U2_n274, B => U2_x_10_6_port, C => U2_n275, D 
                           => U2_x_11_6_port, Q => U2_n520);
   U194 : AOI220 port map( A => U2_n276, B => U2_x_8_6_port, C => U2_n277, D =>
                           U2_x_9_6_port, Q => U2_n521);
   U195 : AOI220 port map( A => U2_n270, B => U2_x_14_6_port, C => U2_n271, D 
                           => U2_x_15_6_port, Q => U2_n518);
   U196 : AOI220 port map( A => U2_n274, B => U2_x_26_7_port, C => U2_n275, D 
                           => U2_x_27_7_port, Q => U2_n364);
   U197 : AOI220 port map( A => U2_n276, B => U2_x_24_7_port, C => U2_n277, D 
                           => U2_x_25_7_port, Q => U2_n365);
   U198 : AOI220 port map( A => U2_n270, B => U2_x_30_7_port, C => U2_n271, D 
                           => U2_x_31_7_port, Q => U2_n362);
   U199 : AOI220 port map( A => U2_n272, B => U2_x_28_6_port, C => U2_n273, D 
                           => U2_x_29_6_port, Q => U2_n385);
   U200 : AOI220 port map( A => U2_n272, B => U2_x_12_6_port, C => U2_n273, D 
                           => U2_x_13_6_port, Q => U2_n519);
   U201 : AOI220 port map( A => U2_n266, B => U2_x_18_7_port, C => U2_n267, D 
                           => U2_x_19_7_port, Q => U2_n360);
   U202 : AOI220 port map( A => U2_n268, B => U2_x_16_7_port, C => U2_n269, D 
                           => U2_x_17_7_port, Q => U2_n361);
   U203 : AOI220 port map( A => U2_n268, B => U2_x_0_7_port, C => U2_n269, D =>
                           U2_x_1_7_port, Q => U2_n371);
   U204 : AOI220 port map( A => U2_n266, B => U2_x_2_7_port, C => U2_n267, D =>
                           U2_x_3_7_port, Q => U2_n370);
   U205 : AOI220 port map( A => U2_n276, B => U2_x_8_7_port, C => U2_n277, D =>
                           U2_x_9_7_port, Q => U2_n375);
   U206 : AOI220 port map( A => U2_n274, B => U2_x_10_7_port, C => U2_n275, D 
                           => U2_x_11_7_port, Q => U2_n374);
   U207 : AOI220 port map( A => U2_n270, B => U2_x_14_7_port, C => U2_n271, D 
                           => U2_x_15_7_port, Q => U2_n372);
   U208 : AOI220 port map( A => U2_n272, B => U2_x_28_7_port, C => U2_n273, D 
                           => U2_x_29_7_port, Q => U2_n363);
   U209 : AOI220 port map( A => U2_n272, B => U2_x_12_7_port, C => U2_n273, D 
                           => U2_x_13_7_port, Q => U2_n373);
   U210 : NAND20 port map( A => n229, B => n121, Q => U6_n43);
   U211 : NAND30 port map( A => U6_n4, B => n19, C => n229, Q => U6_n35);
   U212 : NAND30 port map( A => U6_n2, B => U6_n14, C => U6_n50, Q => U6_n23);
   U213 : OAI210 port map( A => U6_n50, B => U6_n2, C => U6_n23, Q => U6_n31);
   U214 : NAND33 port map( A => U6_n14, B => n30, C => U6_n2, Q => U6_n44);
   U215 : INV3 port map( A => U3_mult_19_FS_1_n27, Q => U3_mult_19_FS_1_n37);
   U216 : INV3 port map( A => n250, Q => n260);
   U217 : INV3 port map( A => n249, Q => n259);
   U218 : INV3 port map( A => n249, Q => n258);
   U219 : INV3 port map( A => n249, Q => n257);
   U220 : INV3 port map( A => n250, Q => n256);
   U221 : INV3 port map( A => U2_n286, Q => n255);
   U222 : INV3 port map( A => n249, Q => n254);
   U223 : INV3 port map( A => n250, Q => n253);
   U224 : INV3 port map( A => n250, Q => n252);
   U225 : INV3 port map( A => n249, Q => n251);
   U226 : INV3 port map( A => Rom_out_7_port, Q => U3_mult_19_n84);
   U227 : NAND22 port map( A => U3_mult_19_A2_7_port, B => U3_mult_19_A1_7_port
                           , Q => U3_mult_19_FS_1_n12);
   U228 : AOI211 port map( A => U3_mult_19_FS_1_n33, B => U3_mult_19_A1_12_port
                           , C => U3_mult_19_FS_1_n32, Q => U3_mult_19_FS_1_n17
                           );
   U229 : INV3 port map( A => U3_mult_19_FS_1_n18, Q => U3_mult_19_FS_1_n32);
   U230 : BUF2 port map( A => U2_n357, Q => n235);
   U231 : IMUX21 port map( A => U3_mult_19_FS_1_n15, B => U3_mult_19_FS_1_n16, 
                           S => U3_mult_19_A2_8_port, Q => U3_mult_19_FS_1_n14)
                           ;
   U232 : XNR21 port map( A => U3_mult_19_A1_8_port, B => U3_mult_19_FS_1_n12, 
                           Q => U3_mult_19_FS_1_n15);
   U233 : INV3 port map( A => U3_mult_19_FS_1_n19, Q => U3_mult_19_FS_1_n33);
   U234 : AOI2111 port map( A => U3_mult_19_FS_1_n20, B => 
                           U3_mult_19_A1_11_port, C => U3_mult_19_FS_1_n34, D 
                           => U3_mult_19_FS_1_n21, Q => U3_mult_19_FS_1_n19);
   U235 : NOR40 port map( A => U3_mult_19_FS_1_n22, B => U3_mult_19_FS_1_n12, C
                           => U3_mult_19_FS_1_n23, D => U3_mult_19_FS_1_n24, Q 
                           => U3_mult_19_FS_1_n21);
   U236 : INV3 port map( A => U3_mult_19_FS_1_n25, Q => U3_mult_19_FS_1_n34);
   U237 : NOR21 port map( A => U3_mult_19_A2_10_port, B => 
                           U3_mult_19_A1_10_port, Q => U3_mult_19_FS_1_n23);
   U238 : NAND22 port map( A => U3_mult_19_A2_9_port, B => U3_mult_19_A1_9_port
                           , Q => U3_mult_19_FS_1_n11);
   U239 : NOR21 port map( A => U3_mult_19_A2_9_port, B => U3_mult_19_A1_9_port,
                           Q => U3_mult_19_FS_1_n22);
   U240 : NAND22 port map( A => U3_mult_19_A2_10_port, B => 
                           U3_mult_19_A1_10_port, Q => U3_mult_19_FS_1_n26);
   U241 : INV3 port map( A => U1_n16, Q => U1_n6);
   U242 : INV3 port map( A => n248, Q => n244);
   U243 : INV3 port map( A => n245, Q => n243);
   U244 : INV3 port map( A => n246, Q => n242);
   U245 : INV3 port map( A => n246, Q => n241);
   U246 : INV3 port map( A => n245, Q => n240);
   U247 : INV3 port map( A => n245, Q => n239);
   U248 : INV3 port map( A => n248, Q => n238);
   U249 : INV3 port map( A => n246, Q => n237);
   U250 : BUF2 port map( A => n250, Q => n261);
   U251 : BUF2 port map( A => n249, Q => n262);
   U252 : XOR21 port map( A => U3_mult_19_SUMB_7_3_port, B => 
                           U3_mult_19_CARRYB_7_2_port, Q => 
                           U3_mult_19_A1_8_port);
   U253 : XOR21 port map( A => U3_mult_19_SUMB_7_2_port, B => 
                           U3_mult_19_CARRYB_7_1_port, Q => 
                           U3_mult_19_A1_7_port);
   U254 : NOR21 port map( A => U2_n278, B => n232, Q => U2_n738);
   U255 : NOR21 port map( A => U2_n278, B => Rom_Address_2_port, Q => U2_n733);
   U256 : INV3 port map( A => U2_n727, Q => U2_n266);
   U257 : INV3 port map( A => U2_n726, Q => U2_n267);
   U258 : INV3 port map( A => U2_n740, Q => U2_n271);
   U259 : NAND22 port map( A => U2_n738, B => U2_n718, Q => U2_n740);
   U260 : NOR21 port map( A => U1_n20, B => n233, Q => U1_n24);
   U261 : NOR21 port map( A => U1_n2, B => n233, Q => U1_n17);
   U262 : AOI211 port map( A => U1_n15, B => U1_n7, C => U1_n24, Q => U1_n31);
   U263 : INV3 port map( A => U2_n736, Q => U2_n274);
   U264 : NAND22 port map( A => U2_n733, B => U2_n717, Q => U2_n736);
   U265 : INV3 port map( A => U2_n735, Q => U2_n275);
   U266 : NAND22 port map( A => U2_n733, B => U2_n718, Q => U2_n735);
   U267 : NAND22 port map( A => U2_n716, B => U2_n718, Q => U2_n356);
   U268 : INV3 port map( A => U1_n37, Q => Rom_out_7_port);
   U269 : INV3 port map( A => U3_mult_19_ab_0_5_port, Q => U3_mult_19_n80);
   U270 : INV3 port map( A => U3_mult_19_ab_0_3_port, Q => U3_mult_19_n78);
   U271 : INV3 port map( A => U3_mult_19_ab_1_4_port, Q => U3_mult_19_n72);
   U272 : INV3 port map( A => U3_mult_19_ab_1_3_port, Q => U3_mult_19_n71);
   U273 : INV3 port map( A => Rom_out_0_port, Q => U3_mult_19_n91);
   U274 : OAI2111 port map( A => U1_n18, B => U1_n4, C => U1_n11, D => U1_n52, 
                           Q => Rom_out_0_port);
   U275 : INV3 port map( A => U1_n24, Q => U1_n4);
   U276 : AOI311 port map( A => U1_n16, B => U1_n7, C => U1_n15, D => U1_n53, Q
                           => U1_n52);
   U277 : XOR21 port map( A => U3_mult_19_SUMB_7_4_port, B => 
                           U3_mult_19_CARRYB_7_3_port, Q => 
                           U3_mult_19_A1_9_port);
   U278 : XOR21 port map( A => U3_mult_19_SUMB_7_5_port, B => 
                           U3_mult_19_CARRYB_7_4_port, Q => 
                           U3_mult_19_A1_10_port);
   U279 : INV3 port map( A => Rom_out_2_port, Q => U3_mult_19_n89);
   U280 : NAND22 port map( A => U1_n41, B => U1_n42, Q => Rom_out_2_port);
   U281 : AOI221 port map( A => U1_n44, B => U1_n2, C => n233, D => U1_n45, Q 
                           => U1_n41);
   U282 : AOI311 port map( A => n232, B => U1_n7, C => U1_n11, D => U1_n43, Q 
                           => U1_n42);
   U283 : NAND22 port map( A => U1_n9, B => U1_n7, Q => U1_n16);
   U284 : NOR21 port map( A => U1_n19, B => U1_n7, Q => U1_n35);
   U285 : NOR21 port map( A => U3_mult_19_n51, B => U3_mult_19_n54, Q => 
                           U3_mult_19_A2_9_port);
   U286 : INV3 port map( A => U3_mult_19_CARRYB_7_2_port, Q => U3_mult_19_n51);
   U287 : INV3 port map( A => U3_mult_19_SUMB_7_3_port, Q => U3_mult_19_n54);
   U288 : NOR31 port map( A => U1_n3, B => U1_n28, C => U1_n35, Q => U1_n53);
   U289 : INV3 port map( A => U1_n25, Q => U1_n3);
   U290 : BUF2 port map( A => U2_n359, Q => n236);
   U291 : INV3 port map( A => U1_n19, Q => U1_n9);
   U292 : INV3 port map( A => U1_n18, Q => U1_n5);
   U293 : XOR21 port map( A => U3_mult_19_SUMB_7_6_port, B => 
                           U3_mult_19_CARRYB_7_5_port, Q => 
                           U3_mult_19_A1_11_port);
   U294 : INV3 port map( A => Mult_out_0_port, Q => U4_add_27_aco_n20);
   U295 : XOR21 port map( A => U3_mult_19_ab_7_7_port, B => 
                           U3_mult_19_CARRYB_7_6_port, Q => 
                           U3_mult_19_A1_12_port);
   U296 : BUF2 port map( A => U2_n286, Q => n250);
   U297 : BUF2 port map( A => U2_n286, Q => n249);
   U298 : BUF2 port map( A => U2_n285, Q => n245);
   U299 : BUF2 port map( A => U2_n285, Q => n248);
   U300 : BUF2 port map( A => U2_n285, Q => n246);
   U301 : BUF2 port map( A => n246, Q => n247);
   U302 : INV3 port map( A => Rom_out_5_port, Q => U3_mult_19_n86);
   U303 : OAI2111 port map( A => U1_n19, B => U1_n20, C => U1_n21, D => U1_n22,
                           Q => Rom_out_5_port);
   U304 : INV3 port map( A => Rom_out_6_port, Q => U3_mult_19_n85);
   U305 : NAND22 port map( A => U1_n13, B => U1_n14, Q => Rom_out_6_port);
   U306 : AOI221 port map( A => U1_n18, B => U1_n2, C => U1_n6, D => 
                           Rom_Address_4_port, Q => U1_n13);
   U307 : AOI221 port map( A => U1_n15, B => U1_n16, C => U1_n17, D => U1_n5, Q
                           => U1_n14);
   U308 : XNR21 port map( A => Rom_Address_4_port, B => n233, Q => U1_n25);
   U309 : NOR21 port map( A => U2_n280, B => n230, Q => U2_n717);
   U310 : NOR21 port map( A => U2_n280, B => U1_n12, Q => U2_n718);
   U311 : NOR21 port map( A => U3_mult_19_n62, B => U3_mult_19_n91, Q => 
                           U3_mult_19_ab_7_0_port);
   U312 : NOR21 port map( A => U3_mult_19_n62, B => U3_mult_19_n90, Q => 
                           U3_mult_19_ab_7_1_port);
   U313 : NOR21 port map( A => n233, B => n231, Q => U2_n724);
   U314 : NOR21 port map( A => U3_mult_19_n62, B => U3_mult_19_n89, Q => 
                           U3_mult_19_ab_7_2_port);
   U315 : NOR21 port map( A => U3_mult_19_n62, B => U3_mult_19_n88, Q => 
                           U3_mult_19_ab_7_3_port);
   U316 : INV3 port map( A => Rom_out_4_port, Q => U3_mult_19_n87);
   U317 : OAI2111 port map( A => U1_n31, B => U1_n32, C => U1_n33, D => U1_n34,
                           Q => Rom_out_4_port);
   U318 : NAND22 port map( A => U1_n35, B => U1_n15, Q => U1_n33);
   U319 : AOI221 port map( A => U1_n28, B => U1_n17, C => U1_n25, D => U1_n32, 
                           Q => U1_n34);
   U320 : INV3 port map( A => U2_n732, Q => U2_n277);
   U321 : NAND22 port map( A => U2_n733, B => U2_n720, Q => U2_n732);
   U322 : INV3 port map( A => Rom_Address_4_port, Q => U1_n2);
   U323 : NOR21 port map( A => U3_mult_19_n91, B => U3_mult_19_n65, Q => 
                           U3_mult_19_ab_4_0_port);
   U324 : NOR21 port map( A => U3_mult_19_n90, B => U3_mult_19_n65, Q => 
                           U3_mult_19_ab_4_1_port);
   U325 : NOR21 port map( A => U3_mult_19_n89, B => U3_mult_19_n65, Q => 
                           U3_mult_19_ab_4_2_port);
   U326 : NOR21 port map( A => U3_mult_19_n88, B => U3_mult_19_n65, Q => 
                           U3_mult_19_ab_4_3_port);
   U327 : NOR21 port map( A => U3_mult_19_n87, B => U3_mult_19_n65, Q => 
                           U3_mult_19_ab_4_4_port);
   U328 : NOR21 port map( A => U3_mult_19_n91, B => U3_mult_19_n64, Q => 
                           U3_mult_19_ab_5_0_port);
   U329 : NOR21 port map( A => U3_mult_19_n90, B => U3_mult_19_n64, Q => 
                           U3_mult_19_ab_5_1_port);
   U330 : NOR21 port map( A => U3_mult_19_n89, B => U3_mult_19_n64, Q => 
                           U3_mult_19_ab_5_2_port);
   U331 : NOR21 port map( A => U3_mult_19_n88, B => U3_mult_19_n64, Q => 
                           U3_mult_19_ab_5_3_port);
   U332 : NOR21 port map( A => U3_mult_19_n91, B => U3_mult_19_n63, Q => 
                           U3_mult_19_ab_6_0_port);
   U333 : NOR21 port map( A => U3_mult_19_n90, B => U3_mult_19_n63, Q => 
                           U3_mult_19_ab_6_1_port);
   U334 : NOR21 port map( A => U3_mult_19_n89, B => U3_mult_19_n63, Q => 
                           U3_mult_19_ab_6_2_port);
   U335 : NOR21 port map( A => U3_mult_19_n88, B => U3_mult_19_n63, Q => 
                           U3_mult_19_ab_6_3_port);
   U336 : NOR21 port map( A => U3_mult_19_n90, B => U3_mult_19_n66, Q => 
                           U3_mult_19_ab_3_1_port);
   U337 : NOR21 port map( A => U3_mult_19_n89, B => U3_mult_19_n66, Q => 
                           U3_mult_19_ab_3_2_port);
   U338 : NOR21 port map( A => U3_mult_19_n88, B => U3_mult_19_n66, Q => 
                           U3_mult_19_ab_3_3_port);
   U339 : NOR21 port map( A => U3_mult_19_n87, B => U3_mult_19_n66, Q => 
                           U3_mult_19_ab_3_4_port);
   U340 : NOR21 port map( A => U3_mult_19_n86, B => U3_mult_19_n66, Q => 
                           U3_mult_19_ab_3_5_port);
   U341 : NOR21 port map( A => U3_mult_19_n90, B => U3_mult_19_n67, Q => 
                           U3_mult_19_ab_2_1_port);
   U342 : XOR21 port map( A => U3_mult_19_ab_0_3_port, B => 
                           U3_mult_19_ab_1_2_port, Q => 
                           U3_mult_19_SUMB_1_2_port);
   U343 : NOR21 port map( A => U3_mult_19_n89, B => U3_mult_19_n67, Q => 
                           U3_mult_19_ab_2_2_port);
   U344 : NOR21 port map( A => U3_mult_19_n78, B => U3_mult_19_n70, Q => 
                           U3_mult_19_CARRYB_1_2_port);
   U345 : XOR21 port map( A => U3_mult_19_ab_0_4_port, B => 
                           U3_mult_19_ab_1_3_port, Q => 
                           U3_mult_19_SUMB_1_3_port);
   U346 : NOR21 port map( A => U3_mult_19_n88, B => U3_mult_19_n67, Q => 
                           U3_mult_19_ab_2_3_port);
   U347 : NOR21 port map( A => U3_mult_19_n79, B => U3_mult_19_n71, Q => 
                           U3_mult_19_CARRYB_1_3_port);
   U348 : XOR21 port map( A => U3_mult_19_ab_0_5_port, B => 
                           U3_mult_19_ab_1_4_port, Q => 
                           U3_mult_19_SUMB_1_4_port);
   U349 : NOR21 port map( A => U3_mult_19_n87, B => U3_mult_19_n67, Q => 
                           U3_mult_19_ab_2_4_port);
   U350 : NOR21 port map( A => U3_mult_19_n80, B => U3_mult_19_n72, Q => 
                           U3_mult_19_CARRYB_1_4_port);
   U351 : XOR21 port map( A => U3_mult_19_ab_0_6_port, B => 
                           U3_mult_19_ab_1_5_port, Q => 
                           U3_mult_19_SUMB_1_5_port);
   U352 : NOR21 port map( A => U3_mult_19_n86, B => U3_mult_19_n67, Q => 
                           U3_mult_19_ab_2_5_port);
   U353 : XOR21 port map( A => U3_mult_19_ab_0_7_port, B => 
                           U3_mult_19_ab_1_6_port, Q => 
                           U3_mult_19_SUMB_1_6_port);
   U354 : NOR21 port map( A => U3_mult_19_n87, B => U3_mult_19_n75, Q => 
                           U3_mult_19_ab_1_4_port);
   U355 : NOR21 port map( A => U3_mult_19_n86, B => U3_mult_19_n75, Q => 
                           U3_mult_19_ab_1_5_port);
   U356 : NOR21 port map( A => U3_mult_19_n85, B => U3_mult_19_n75, Q => 
                           U3_mult_19_ab_1_6_port);
   U357 : NOR21 port map( A => U3_mult_19_n86, B => U3_mult_19_n83, Q => 
                           U3_mult_19_ab_0_5_port);
   U358 : NOR21 port map( A => U3_mult_19_n85, B => U3_mult_19_n83, Q => 
                           U3_mult_19_ab_0_6_port);
   U359 : NOR21 port map( A => U3_mult_19_n84, B => U3_mult_19_n83, Q => 
                           U3_mult_19_ab_0_7_port);
   U360 : INV3 port map( A => U2_n739, Q => U2_n272);
   U361 : NAND22 port map( A => U2_n738, B => U2_n719, Q => U2_n739);
   U362 : NOR21 port map( A => U3_mult_19_n84, B => U3_mult_19_n67, Q => 
                           U3_mult_19_ab_2_7_port);
   U363 : NOR21 port map( A => U3_mult_19_n85, B => U3_mult_19_n66, Q => 
                           U3_mult_19_ab_3_6_port);
   U364 : NOR21 port map( A => U3_mult_19_n86, B => U3_mult_19_n65, Q => 
                           U3_mult_19_ab_4_5_port);
   U365 : NOR21 port map( A => U3_mult_19_n84, B => U3_mult_19_n66, Q => 
                           U3_mult_19_ab_3_7_port);
   U366 : NOR21 port map( A => U3_mult_19_n85, B => U3_mult_19_n65, Q => 
                           U3_mult_19_ab_4_6_port);
   U367 : NOR21 port map( A => U3_mult_19_n87, B => U3_mult_19_n64, Q => 
                           U3_mult_19_ab_5_4_port);
   U368 : NOR21 port map( A => U3_mult_19_n86, B => U3_mult_19_n64, Q => 
                           U3_mult_19_ab_5_5_port);
   U369 : NOR21 port map( A => U3_mult_19_n87, B => U3_mult_19_n63, Q => 
                           U3_mult_19_ab_6_4_port);
   U370 : INV3 port map( A => n232, Q => n233);
   U371 : NOR21 port map( A => U3_mult_19_n85, B => U3_mult_19_n67, Q => 
                           U3_mult_19_ab_2_6_port);
   U372 : INV3 port map( A => Rom_out_3_port, Q => U3_mult_19_n88);
   U373 : AOI2111 port map( A => U1_n9, B => U1_n20, C => U1_n38, D => U1_n39, 
                           Q => U1_n36);
   U374 : XNR21 port map( A => U2_n280, B => n233, Q => U1_n38);
   U375 : NOR21 port map( A => U3_mult_19_n62, B => U3_mult_19_n87, Q => 
                           U3_mult_19_ab_7_4_port);
   U376 : NOR21 port map( A => U3_mult_19_n62, B => U3_mult_19_n86, Q => 
                           U3_mult_19_ab_7_5_port);
   U377 : NOR21 port map( A => n232, B => Rom_Address_4_port, Q => U1_n15);
   U378 : OAI2111 port map( A => U1_n7, B => U1_n32, C => U1_n20, D => U1_n46, 
                           Q => U1_n45);
   U379 : NAND22 port map( A => Rom_Address_4_port, B => U1_n12, Q => U1_n46);
   U380 : NOR21 port map( A => U1_n40, B => U1_n7, Q => U1_n18);
   U381 : NAND22 port map( A => U1_n12, B => U2_n280, Q => U1_n19);
   U382 : NOR21 port map( A => U3_mult_19_n91, B => U3_mult_19_n66, Q => 
                           U3_mult_19_ab_3_0_port);
   U383 : NOR21 port map( A => U3_mult_19_n91, B => U3_mult_19_n67, Q => 
                           U3_mult_19_ab_2_0_port);
   U384 : XOR21 port map( A => U3_mult_19_ab_0_2_port, B => 
                           U3_mult_19_ab_1_1_port, Q => 
                           U3_mult_19_SUMB_1_1_port);
   U385 : AOI211 port map( A => U1_n29, B => U1_n30, C => U1_n7, Q => U1_n27);
   U386 : INV3 port map( A => Rom_out_1_port, Q => U3_mult_19_n90);
   U387 : AOI221 port map( A => n233, B => U1_n50, C => U1_n6, D => U1_n17, Q 
                           => U1_n49);
   U388 : NOR21 port map( A => U3_mult_19_n84, B => U3_mult_19_n65, Q => 
                           U3_mult_19_ab_4_7_port);
   U389 : NOR21 port map( A => U3_mult_19_n85, B => U3_mult_19_n64, Q => 
                           U3_mult_19_ab_5_6_port);
   U390 : NOR21 port map( A => U3_mult_19_n86, B => U3_mult_19_n63, Q => 
                           U3_mult_19_ab_6_5_port);
   U391 : NOR21 port map( A => U3_mult_19_n84, B => U3_mult_19_n64, Q => 
                           U3_mult_19_ab_5_7_port);
   U392 : NOR21 port map( A => U3_mult_19_n85, B => U3_mult_19_n63, Q => 
                           U3_mult_19_ab_6_6_port);
   U393 : INV3 port map( A => U1_n32, Q => U1_n11);
   U394 : NOR21 port map( A => U1_n40, B => U1_n20, Q => U1_n39);
   U395 : NOR21 port map( A => U3_mult_19_n84, B => U3_mult_19_n63, Q => 
                           U3_mult_19_ab_6_7_port);
   U396 : NOR21 port map( A => U3_mult_19_n62, B => U3_mult_19_n85, Q => 
                           U3_mult_19_ab_7_6_port);
   U397 : NOR21 port map( A => U3_mult_19_n62, B => U3_mult_19_n84, Q => 
                           U3_mult_19_ab_7_7_port);
   U398 : NOR21 port map( A => RESET, B => U4_n42, Q => U4_N28_port);
   U399 : INV3 port map( A => U4_N7, Q => U4_n42);
   U400 : NOR21 port map( A => RESET, B => U2_n285, Q => U2_n286);
   U401 : INV3 port map( A => U6_n28, Q => U6_n7);
   U402 : NOR22 port map( A => U5_n11, B => RESET, Q => U5_n3);
   U403 : INV3 port map( A => U5_n11, Q => U5_n1);
   U404 : INV3 port map( A => U8_n5, Q => U8_n1);
   U405 : NOR21 port map( A => n230, B => n229, Q => U2_n719);
   U406 : NOR21 port map( A => U1_n12, B => n229, Q => U2_n720);
   U407 : INV3 port map( A => U6_n29, Q => Rom_Address_4_port);
   U408 : NOR40 port map( A => U2_n712, B => U2_n713, C => U2_n714, D => 
                           U2_n715, Q => U2_n700);
   U409 : NOR40 port map( A => U2_n702, B => U2_n703, C => U2_n704, D => 
                           U2_n705, Q => U2_n701);
   U410 : INV3 port map( A => Delay_Line_out_2_port, Q => U3_mult_19_n67);
   U411 : NOR40 port map( A => U2_n668, B => U2_n669, C => U2_n670, D => 
                           U2_n671, Q => U2_n656);
   U412 : NOR40 port map( A => U2_n658, B => U2_n659, C => U2_n660, D => 
                           U2_n661, Q => U2_n657);
   U413 : NOR40 port map( A => U2_n690, B => U2_n691, C => U2_n692, D => 
                           U2_n693, Q => U2_n678);
   U414 : NOR40 port map( A => U2_n680, B => U2_n681, C => U2_n682, D => 
                           U2_n683, Q => U2_n679);
   U415 : INV3 port map( A => Delay_Line_out_3_port, Q => U3_mult_19_n66);
   U416 : NOR40 port map( A => U2_n646, B => U2_n647, C => U2_n648, D => 
                           U2_n649, Q => U2_n634);
   U417 : NOR40 port map( A => U2_n636, B => U2_n637, C => U2_n638, D => 
                           U2_n639, Q => U2_n635);
   U418 : NOR21 port map( A => RESET, B => n224, Q => U4_N46);
   U419 : INV3 port map( A => U6_n44, Q => U6_n11);
   U420 : INV3 port map( A => Rom_Address_2_port, Q => n232);
   U421 : NOR21 port map( A => n19, B => U6_n44, Q => Rom_Address_2_port);
   U422 : BUF2 port map( A => Rom_Address_3_port, Q => n231);
   U423 : NOR21 port map( A => n31, B => U6_n44, Q => Rom_Address_3_port);
   U424 : NOR21 port map( A => U4_add_27_aco_n14, B => 
                           U4_mult_add_27_aco_PROD_not_18_port, Q => 
                           U4_add_27_aco_carry_19_port);
   U425 : INV3 port map( A => U4_add_27_aco_carry_18_port, Q => 
                           U4_add_27_aco_n14);
   U426 : NOR21 port map( A => U4_add_27_aco_n18, B => 
                           U4_mult_add_27_aco_PROD_not_16_port, Q => 
                           U4_add_27_aco_carry_17_port);
   U427 : NOR40 port map( A => U2_n624, B => U2_n625, C => U2_n626, D => 
                           U2_n627, Q => U2_n612);
   U428 : NOR40 port map( A => U2_n614, B => U2_n615, C => U2_n616, D => 
                           U2_n617, Q => U2_n613);
   U429 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_1_port, Q => U4_N49);
   U430 : NOR21 port map( A => U4_add_27_aco_n20, B => 
                           U4_mult_add_27_aco_PROD_not_0_port, Q => 
                           U4_add_27_aco_carry_1_port);
   U431 : XOR21 port map( A => U3_mult_19_ab_0_1_port, B => 
                           U3_mult_19_ab_1_0_port, Q => Mult_out_1_port);
   U432 : NOR21 port map( A => RESET, B => U4_n29, Q => U4_N41_port);
   U433 : INV3 port map( A => U4_N20, Q => U4_n29);
   U434 : NOR21 port map( A => RESET, B => U4_n28, Q => U4_N42_port);
   U435 : INV3 port map( A => U4_N21, Q => U4_n28);
   U436 : NOR40 port map( A => U2_n602, B => U2_n603, C => U2_n604, D => 
                           U2_n605, Q => U2_n522);
   U437 : NOR40 port map( A => U2_n592, B => U2_n593, C => U2_n594, D => 
                           U2_n595, Q => U2_n523);
   U438 : INV3 port map( A => Delay_Line_out_6_port, Q => U3_mult_19_n63);
   U439 : NOR40 port map( A => U2_n388, B => U2_n389, C => U2_n390, D => 
                           U2_n391, Q => U2_n376);
   U440 : NOR40 port map( A => U2_n378, B => U2_n379, C => U2_n380, D => 
                           U2_n381, Q => U2_n377);
   U441 : NOR21 port map( A => RESET, B => U4_n30, Q => U4_N40_port);
   U442 : INV3 port map( A => U4_N19, Q => U4_n30);
   U443 : NOR21 port map( A => RESET, B => U4_n31, Q => U4_N39_port);
   U444 : INV3 port map( A => U4_N18, Q => U4_n31);
   U445 : NOR21 port map( A => RESET, B => U4_n32, Q => U4_N38_port);
   U446 : INV3 port map( A => U4_N17, Q => U4_n32);
   U447 : NOR40 port map( A => U2_n366, B => U2_n367, C => U2_n368, D => 
                           U2_n369, Q => U2_n350);
   U448 : NOR40 port map( A => U2_n352, B => U2_n353, C => U2_n354, D => 
                           U2_n355, Q => U2_n351);
   U449 : NOR21 port map( A => RESET, B => U4_n33, Q => U4_N37_port);
   U450 : INV3 port map( A => U4_N16, Q => U4_n33);
   U451 : BUF2 port map( A => U6_n24, Q => n234);
   U452 : NOR21 port map( A => RESET, B => U4_n35, Q => U4_N35_port);
   U453 : INV3 port map( A => U4_N14, Q => U4_n35);
   U454 : NOR21 port map( A => RESET, B => U4_n34, Q => U4_N36_port);
   U455 : INV3 port map( A => U4_N15, Q => U4_n34);
   U456 : NOR21 port map( A => RESET, B => U4_n36, Q => U4_N34_port);
   U457 : INV3 port map( A => U4_N13, Q => U4_n36);
   U458 : NOR21 port map( A => RESET, B => U4_n37, Q => U4_N33_port);
   U459 : INV3 port map( A => U4_N12, Q => U4_n37);
   U460 : NOR21 port map( A => RESET, B => U4_n39, Q => U4_N31_port);
   U461 : INV3 port map( A => U4_N10, Q => U4_n39);
   U462 : NOR21 port map( A => RESET, B => U4_n38, Q => U4_N32_port);
   U463 : INV3 port map( A => U4_N11, Q => U4_n38);
   U464 : NOR21 port map( A => RESET, B => U4_n40, Q => U4_N30_port);
   U465 : INV3 port map( A => U4_N9, Q => U4_n40);
   U466 : NOR21 port map( A => RESET, B => U4_n41, Q => U4_N29_port);
   U467 : INV3 port map( A => U4_N8, Q => U4_n41);
   U468 : INV3 port map( A => ack_F2ADC, Q => U6_n16);
   U469 : NOR21 port map( A => RESET, B => Delay_Line_sample_shift, Q => 
                           U2_n285);
   U470 : OAI2111 port map( A => U6_n27, B => U1_n7, C => U6_n32, D => U6_n34, 
                           Q => U6_n40);
   U471 : NAND31 port map( A => U6_n11, B => n31, C => U6_n27, Q => U6_n32);
   U472 : NAND31 port map( A => U6_n16, B => U6_n28, C => U6_n46, Q => U6_n37);
   U473 : AOI211 port map( A => U6_n11, B => n121, C => U6_n31, Q => U6_n46);
   U474 : NOR21 port map( A => Buff_OE, B => U6_n8, Q => U6_n28);
   U475 : INV3 port map( A => U6_n34, Q => U6_n8);
   U476 : NOR22 port map( A => U9_n11, B => RESET, Q => U9_n3);
   U477 : INV3 port map( A => U9_n11, Q => U9_n1);
   U478 : NOR21 port map( A => Buff_OE, B => RESET, Q => U5_n11);
   U479 : INV3 port map( A => U6_n27, Q => U6_n13);
   U480 : NAND22 port map( A => req_F2DAC, B => n263, Q => U8_n5);
   U481 : INV3 port map( A => U6_n23, Q => req_F2DAC);
   U482 : INV3 port map( A => U7_n12, Q => req_ADC2F);
   U483 : NOR21 port map( A => req_ADC2F, B => U7_n1, Q => U7_n14);
   U484 : INV3 port map( A => ADC_Rdb_port, Q => U7_n1);
   U485 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_15_port, Q => U4_N63)
                           ;
   U486 : NAND22 port map( A => Accu_out_15_port, B => U6_n24, Q => 
                           U4_mult_add_27_aco_PROD_not_15_port);
   U487 : NAND41 port map( A => U2_n708, B => U2_n709, C => U2_n710, D => 
                           U2_n711, Q => U2_n702);
   U488 : AOI221 port map( A => U2_n274, B => U2_x_26_0_port, C => U2_n275, D 
                           => U2_x_27_0_port, Q => U2_n710);
   U489 : AOI221 port map( A => U2_n276, B => U2_x_24_0_port, C => U2_n277, D 
                           => U2_x_25_0_port, Q => U2_n711);
   U490 : AOI221 port map( A => U2_n270, B => U2_x_30_0_port, C => U2_n271, D 
                           => U2_x_31_0_port, Q => U2_n708);
   U491 : NAND41 port map( A => U2_n728, B => U2_n729, C => U2_n730, D => 
                           U2_n731, Q => U2_n712);
   U492 : NAND41 port map( A => U2_n664, B => U2_n665, C => U2_n666, D => 
                           U2_n667, Q => U2_n658);
   U493 : NAND41 port map( A => U2_n674, B => U2_n675, C => U2_n676, D => 
                           U2_n677, Q => U2_n668);
   U494 : NAND41 port map( A => U2_n686, B => U2_n687, C => U2_n688, D => 
                           U2_n689, Q => U2_n680);
   U495 : AOI221 port map( A => U2_n274, B => U2_x_26_1_port, C => U2_n275, D 
                           => U2_x_27_1_port, Q => U2_n688);
   U496 : AOI221 port map( A => U2_n276, B => U2_x_24_1_port, C => U2_n277, D 
                           => U2_x_25_1_port, Q => U2_n689);
   U497 : AOI221 port map( A => U2_n270, B => U2_x_30_1_port, C => U2_n271, D 
                           => U2_x_31_1_port, Q => U2_n686);
   U498 : NAND41 port map( A => U2_n696, B => U2_n697, C => U2_n698, D => 
                           U2_n699, Q => U2_n690);
   U499 : NAND41 port map( A => U2_n642, B => U2_n643, C => U2_n644, D => 
                           U2_n645, Q => U2_n636);
   U500 : NAND22 port map( A => U6_n48, B => U6_n11, Q => U6_n29);
   U501 : AOI221 port map( A => U2_n272, B => U2_x_28_0_port, C => U2_n273, D 
                           => U2_x_29_0_port, Q => U2_n709);
   U502 : AOI221 port map( A => U2_n272, B => U2_x_28_1_port, C => U2_n273, D 
                           => U2_x_29_1_port, Q => U2_n687);
   U503 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_14_port, Q => U4_N62)
                           ;
   U504 : NAND22 port map( A => Accu_out_14_port, B => n234, Q => 
                           U4_mult_add_27_aco_PROD_not_14_port);
   U505 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_10_port, Q => U4_N58)
                           ;
   U506 : NAND22 port map( A => U4_Accu_out_10_port, B => n234, Q => 
                           U4_mult_add_27_aco_PROD_not_10_port);
   U507 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_8_port, Q => U4_N56);
   U508 : NAND22 port map( A => U4_Accu_out_8_port, B => U6_n24, Q => 
                           U4_mult_add_27_aco_PROD_not_8_port);
   U509 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_12_port, Q => U4_N60)
                           ;
   U510 : NAND22 port map( A => Accu_out_12_port, B => n234, Q => 
                           U4_mult_add_27_aco_PROD_not_12_port);
   U511 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_9_port, Q => U4_N57);
   U512 : NAND22 port map( A => n234, B => U4_Accu_out_9_port, Q => 
                           U4_mult_add_27_aco_PROD_not_9_port);
   U513 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_11_port, Q => U4_N59)
                           ;
   U514 : XNR21 port map( A => U3_mult_19_FS_1_n9, B => U3_mult_19_FS_1_n10, Q 
                           => Mult_out_11_port);
   U515 : NAND22 port map( A => U4_Accu_out_11_port, B => U6_n24, Q => 
                           U4_mult_add_27_aco_PROD_not_11_port);
   U516 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_6_port, Q => U4_N54);
   U517 : NAND22 port map( A => U4_Accu_out_6_port, B => n234, Q => 
                           U4_mult_add_27_aco_PROD_not_6_port);
   U518 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_7_port, Q => U4_N55);
   U519 : NAND22 port map( A => U4_Accu_out_7_port, B => n234, Q => 
                           U4_mult_add_27_aco_PROD_not_7_port);
   U520 : NAND22 port map( A => U2_n706, B => U2_n707, Q => U2_n703);
   U521 : AOI221 port map( A => U2_n266, B => U2_x_18_0_port, C => U2_n267, D 
                           => U2_x_19_0_port, Q => U2_n706);
   U522 : AOI221 port map( A => U2_n268, B => U2_x_16_0_port, C => U2_n269, D 
                           => U2_x_17_0_port, Q => U2_n707);
   U523 : NAND22 port map( A => U2_n721, B => U2_n722, Q => U2_n713);
   U524 : AOI221 port map( A => U2_n266, B => U2_x_2_0_port, C => U2_n267, D =>
                           U2_x_3_0_port, Q => U2_n721);
   U525 : NAND22 port map( A => U2_n662, B => U2_n663, Q => U2_n659);
   U526 : NAND22 port map( A => U2_n672, B => U2_n673, Q => U2_n669);
   U527 : NAND22 port map( A => U2_n684, B => U2_n685, Q => U2_n681);
   U528 : AOI221 port map( A => U2_n266, B => U2_x_18_1_port, C => U2_n267, D 
                           => U2_x_19_1_port, Q => U2_n684);
   U529 : AOI221 port map( A => U2_n268, B => U2_x_16_1_port, C => U2_n269, D 
                           => U2_x_17_1_port, Q => U2_n685);
   U530 : NAND22 port map( A => U2_n694, B => U2_n695, Q => U2_n691);
   U531 : AOI221 port map( A => U2_n266, B => U2_x_2_1_port, C => U2_n267, D =>
                           U2_x_3_1_port, Q => U2_n694);
   U532 : NAND41 port map( A => U2_n652, B => U2_n653, C => U2_n654, D => 
                           U2_n655, Q => U2_n646);
   U533 : NAND41 port map( A => U2_n620, B => U2_n621, C => U2_n622, D => 
                           U2_n623, Q => U2_n614);
   U534 : NAND41 port map( A => U2_n630, B => U2_n631, C => U2_n632, D => 
                           U2_n633, Q => U2_n624);
   U535 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_2_port, Q => U4_N50);
   U536 : NAND22 port map( A => U4_Accu_out_2_port, B => n234, Q => 
                           U4_mult_add_27_aco_PROD_not_2_port);
   U537 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_3_port, Q => U4_N51);
   U538 : NAND22 port map( A => U4_Accu_out_3_port, B => n234, Q => 
                           U4_mult_add_27_aco_PROD_not_3_port);
   U539 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_4_port, Q => U4_N52);
   U540 : NAND22 port map( A => U4_Accu_out_4_port, B => n234, Q => 
                           U4_mult_add_27_aco_PROD_not_4_port);
   U541 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_5_port, Q => U4_N53);
   U542 : NAND22 port map( A => U4_Accu_out_5_port, B => n234, Q => 
                           U4_mult_add_27_aco_PROD_not_5_port);
   U543 : NAND22 port map( A => U2_n640, B => U2_n641, Q => U2_n637);
   U544 : NAND22 port map( A => U2_n650, B => U2_n651, Q => U2_n647);
   U545 : NAND22 port map( A => U2_n618, B => U2_n619, Q => U2_n615);
   U546 : NAND22 port map( A => U2_n628, B => U2_n629, Q => U2_n625);
   U547 : NAND41 port map( A => U2_n598, B => U2_n599, C => U2_n600, D => 
                           U2_n601, Q => U2_n592);
   U548 : NAND41 port map( A => U2_n608, B => U2_n609, C => U2_n610, D => 
                           U2_n611, Q => U2_n602);
   U549 : NAND41 port map( A => U2_n384, B => U2_n385, C => U2_n386, D => 
                           U2_n387, Q => U2_n378);
   U550 : NAND41 port map( A => U2_n518, B => U2_n519, C => U2_n520, D => 
                           U2_n521, Q => U2_n388);
   U551 : NAND22 port map( A => U2_n596, B => U2_n597, Q => U2_n593);
   U552 : NAND22 port map( A => U2_n606, B => U2_n607, Q => U2_n603);
   U553 : NAND22 port map( A => U2_n382, B => U2_n383, Q => U2_n379);
   U554 : NAND22 port map( A => U2_n516, B => U2_n517, Q => U2_n389);
   U555 : NAND41 port map( A => U2_n362, B => U2_n363, C => U2_n364, D => 
                           U2_n365, Q => U2_n352);
   U556 : NAND41 port map( A => U2_n372, B => U2_n373, C => U2_n374, D => 
                           U2_n375, Q => U2_n366);
   U557 : NAND22 port map( A => U2_n360, B => U2_n361, Q => U2_n353);
   U558 : NAND22 port map( A => U2_n370, B => U2_n371, Q => U2_n367);
   U559 : NOR21 port map( A => U6_n14, B => U6_n50, Q => ack_F2ADC);
   U560 : NAND22 port map( A => U4_Accu_out_1_port, B => n234, Q => 
                           U4_mult_add_27_aco_PROD_not_1_port);
   U561 : NAND22 port map( A => U4_Accu_out_0_port, B => U6_n24, Q => 
                           U4_mult_add_27_aco_PROD_not_0_port);
   U562 : NAND22 port map( A => U6_n2, B => ack_F2ADC, Q => U6_n24);
   U563 : NAND31 port map( A => U6_n47, B => U6_n27, C => Rom_Address_4_port, Q
                           => U6_n34);
   U564 : OAI2111 port map( A => U1_n12, B => n223, C => U6_n34, D => U6_n43, Q
                           => U6_n38);
   U565 : INV3 port map( A => U2_n287, Q => U2_n3);
   U566 : AOI221 port map( A => n248, B => U2_x_1_6_port, C => n250, D => 
                           U2_x_0_6_port, Q => U2_n287);
   U567 : INV3 port map( A => U2_n288, Q => U2_n5);
   U568 : AOI221 port map( A => n248, B => U2_x_1_5_port, C => n261, D => 
                           U2_x_0_5_port, Q => U2_n288);
   U569 : NAND31 port map( A => U6_n35, B => U6_n34, C => U6_n36, Q => U6_n39);
   U570 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_16_port, Q => U4_N64)
                           ;
   U571 : NAND22 port map( A => Accu_out_16_port, B => n234, Q => 
                           U4_mult_add_27_aco_PROD_not_16_port);
   U572 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_17_port, Q => U4_N65)
                           ;
   U573 : NAND22 port map( A => Accu_out_17_port, B => U6_n24, Q => 
                           U4_mult_add_27_aco_PROD_not_17_port);
   U574 : INV3 port map( A => U4_mult_add_27_aco_PROD_not_18_port, Q => U4_N66)
                           ;
   U575 : NAND22 port map( A => Accu_out_18_port, B => n234, Q => 
                           U4_mult_add_27_aco_PROD_not_18_port);
   U576 : INV3 port map( A => U2_n349, Q => U2_n2);
   U577 : AOI221 port map( A => U2_x_0_7_port, B => U2_n285, C => n261, D => 
                           Filter_In_mem_7_port, Q => U2_n349);
   U578 : INV3 port map( A => U2_n302, Q => U2_n25);
   U579 : AOI221 port map( A => n246, B => U2_x_3_7_port, C => U2_n286, D => 
                           U2_x_2_7_port, Q => U2_n302);
   U580 : INV3 port map( A => U2_n303, Q => U2_n26);
   U581 : AOI221 port map( A => n248, B => U2_x_3_6_port, C => n262, D => 
                           U2_x_2_6_port, Q => U2_n303);
   U582 : INV3 port map( A => U2_n304, Q => U2_n27);
   U583 : AOI221 port map( A => n248, B => U2_x_3_5_port, C => n261, D => 
                           U2_x_2_5_port, Q => U2_n304);
   U584 : INV3 port map( A => U2_n305, Q => U2_n28);
   U585 : AOI221 port map( A => n247, B => U2_x_3_4_port, C => U2_n286, D => 
                           U2_x_2_4_port, Q => U2_n305);
   U586 : INV3 port map( A => U2_n306, Q => U2_n29);
   U587 : AOI221 port map( A => n246, B => U2_x_3_3_port, C => U2_n286, D => 
                           U2_x_2_3_port, Q => U2_n306);
   U588 : INV3 port map( A => U2_n307, Q => U2_n30);
   U589 : AOI221 port map( A => n245, B => U2_x_3_2_port, C => n261, D => 
                           U2_x_2_2_port, Q => U2_n307);
   U590 : INV3 port map( A => U2_n308, Q => U2_n31);
   U591 : AOI221 port map( A => n246, B => U2_x_3_1_port, C => n250, D => 
                           U2_x_2_1_port, Q => U2_n308);
   U592 : INV3 port map( A => U2_n309, Q => U2_n32);
   U593 : AOI221 port map( A => n246, B => U2_x_3_0_port, C => n262, D => 
                           U2_x_2_0_port, Q => U2_n309);
   U594 : INV3 port map( A => U2_n348, Q => U2_n4);
   U595 : AOI221 port map( A => n246, B => U2_x_0_6_port, C => n262, D => 
                           Filter_In_mem_6_port, Q => U2_n348);
   U596 : INV3 port map( A => U2_n347, Q => U2_n6);
   U597 : AOI221 port map( A => n248, B => U2_x_0_5_port, C => n249, D => 
                           Filter_In_mem_5_port, Q => U2_n347);
   U598 : INV3 port map( A => U2_n346, Q => U2_n8);
   U599 : AOI221 port map( A => n246, B => U2_x_0_4_port, C => n262, D => 
                           Filter_In_mem_4_port, Q => U2_n346);
   U600 : INV3 port map( A => U2_n345, Q => U2_n10);
   U601 : AOI221 port map( A => n247, B => U2_x_0_3_port, C => n249, D => 
                           Filter_In_mem_3_port, Q => U2_n345);
   U602 : INV3 port map( A => U2_n344, Q => U2_n12);
   U603 : AOI221 port map( A => n247, B => U2_x_0_2_port, C => n261, D => 
                           Filter_In_mem_2_port, Q => U2_n344);
   U604 : INV3 port map( A => U2_n343, Q => U2_n14);
   U605 : AOI221 port map( A => n246, B => U2_x_0_1_port, C => n261, D => 
                           Filter_In_mem_1_port, Q => U2_n343);
   U606 : INV3 port map( A => U2_n342, Q => U2_n16);
   U607 : AOI221 port map( A => n245, B => U2_x_0_0_port, C => n261, D => 
                           Filter_In_mem_0_port, Q => U2_n342);
   U608 : INV3 port map( A => U2_n284, Q => U2_n1);
   U609 : AOI221 port map( A => n247, B => U2_x_1_7_port, C => n262, D => 
                           U2_x_0_7_port, Q => U2_n284);
   U610 : INV3 port map( A => U2_n289, Q => U2_n7);
   U611 : AOI221 port map( A => n247, B => U2_x_1_4_port, C => U2_n286, D => 
                           U2_x_0_4_port, Q => U2_n289);
   U612 : INV3 port map( A => U2_n290, Q => U2_n9);
   U613 : AOI221 port map( A => n245, B => U2_x_1_3_port, C => n250, D => 
                           U2_x_0_3_port, Q => U2_n290);
   U614 : INV3 port map( A => U2_n291, Q => U2_n11);
   U615 : AOI221 port map( A => n246, B => U2_x_1_2_port, C => n250, D => 
                           U2_x_0_2_port, Q => U2_n291);
   U616 : INV3 port map( A => U2_n292, Q => U2_n13);
   U617 : AOI221 port map( A => n248, B => U2_x_1_1_port, C => n262, D => 
                           U2_x_0_1_port, Q => U2_n292);
   U618 : INV3 port map( A => U2_n293, Q => U2_n15);
   U619 : AOI221 port map( A => n245, B => U2_x_1_0_port, C => n249, D => 
                           U2_x_0_0_port, Q => U2_n293);
   U620 : INV3 port map( A => U2_n294, Q => U2_n17);
   U621 : AOI221 port map( A => n245, B => U2_x_2_7_port, C => n262, D => 
                           U2_x_1_7_port, Q => U2_n294);
   U622 : INV3 port map( A => U2_n295, Q => U2_n18);
   U623 : AOI221 port map( A => n245, B => U2_x_2_6_port, C => n249, D => 
                           U2_x_1_6_port, Q => U2_n295);
   U624 : INV3 port map( A => U2_n296, Q => U2_n19);
   U625 : AOI221 port map( A => n245, B => U2_x_2_5_port, C => n250, D => 
                           U2_x_1_5_port, Q => U2_n296);
   U626 : INV3 port map( A => U2_n297, Q => U2_n20);
   U627 : AOI221 port map( A => n245, B => U2_x_2_4_port, C => n262, D => 
                           U2_x_1_4_port, Q => U2_n297);
   U628 : INV3 port map( A => U2_n298, Q => U2_n21);
   U629 : AOI221 port map( A => n245, B => U2_x_2_3_port, C => n262, D => 
                           U2_x_1_3_port, Q => U2_n298);
   U630 : INV3 port map( A => U2_n299, Q => U2_n22);
   U631 : AOI221 port map( A => n245, B => U2_x_2_2_port, C => n262, D => 
                           U2_x_1_2_port, Q => U2_n299);
   U632 : INV3 port map( A => U2_n300, Q => U2_n23);
   U633 : AOI221 port map( A => n245, B => U2_x_2_1_port, C => n261, D => 
                           U2_x_1_1_port, Q => U2_n300);
   U634 : INV3 port map( A => U2_n301, Q => U2_n24);
   U635 : AOI221 port map( A => n245, B => U2_x_2_0_port, C => n250, D => 
                           U2_x_1_0_port, Q => U2_n301);
   U636 : INV3 port map( A => U2_n318, Q => U2_n226);
   U637 : AOI221 port map( A => n247, B => U2_x_28_7_port, C => U2_n286, D => 
                           U2_x_27_7_port, Q => U2_n318);
   U638 : INV3 port map( A => U2_n319, Q => U2_n228);
   U639 : AOI221 port map( A => n247, B => U2_x_28_6_port, C => n250, D => 
                           U2_x_27_6_port, Q => U2_n319);
   U640 : INV3 port map( A => U2_n320, Q => U2_n230);
   U641 : AOI221 port map( A => n247, B => U2_x_28_5_port, C => n249, D => 
                           U2_x_27_5_port, Q => U2_n320);
   U642 : INV3 port map( A => U2_n321, Q => U2_n232);
   U643 : AOI221 port map( A => U2_n285, B => U2_x_28_4_port, C => n261, D => 
                           U2_x_27_4_port, Q => U2_n321);
   U644 : INV3 port map( A => U2_n322, Q => U2_n234);
   U645 : AOI221 port map( A => U2_n285, B => U2_x_28_3_port, C => n249, D => 
                           U2_x_27_3_port, Q => U2_n322);
   U646 : INV3 port map( A => U2_n323, Q => U2_n236);
   U647 : AOI221 port map( A => U2_n285, B => U2_x_28_2_port, C => n262, D => 
                           U2_x_27_2_port, Q => U2_n323);
   U648 : INV3 port map( A => U2_n324, Q => U2_n238);
   U649 : AOI221 port map( A => n247, B => U2_x_28_1_port, C => n249, D => 
                           U2_x_27_1_port, Q => U2_n324);
   U650 : INV3 port map( A => U2_n325, Q => U2_n240);
   U651 : AOI221 port map( A => n247, B => U2_x_28_0_port, C => n261, D => 
                           U2_x_27_0_port, Q => U2_n325);
   U652 : INV3 port map( A => U2_n326, Q => U2_n241);
   U653 : AOI221 port map( A => U2_n285, B => U2_x_29_7_port, C => n249, D => 
                           U2_x_28_7_port, Q => U2_n326);
   U654 : INV3 port map( A => U2_n327, Q => U2_n242);
   U655 : AOI221 port map( A => n247, B => U2_x_29_6_port, C => n249, D => 
                           U2_x_28_6_port, Q => U2_n327);
   U656 : INV3 port map( A => U2_n328, Q => U2_n243);
   U657 : AOI221 port map( A => n248, B => U2_x_29_5_port, C => n261, D => 
                           U2_x_28_5_port, Q => U2_n328);
   U658 : INV3 port map( A => U2_n329, Q => U2_n244);
   U659 : AOI221 port map( A => n248, B => U2_x_29_4_port, C => n261, D => 
                           U2_x_28_4_port, Q => U2_n329);
   U660 : INV3 port map( A => U2_n330, Q => U2_n245);
   U661 : AOI221 port map( A => n245, B => U2_x_29_3_port, C => U2_n286, D => 
                           U2_x_28_3_port, Q => U2_n330);
   U662 : INV3 port map( A => U2_n331, Q => U2_n246);
   U663 : AOI221 port map( A => n247, B => U2_x_29_2_port, C => n250, D => 
                           U2_x_28_2_port, Q => U2_n331);
   U664 : INV3 port map( A => U2_n332, Q => U2_n247);
   U665 : AOI221 port map( A => n247, B => U2_x_29_1_port, C => n261, D => 
                           U2_x_28_1_port, Q => U2_n332);
   U666 : INV3 port map( A => U2_n333, Q => U2_n248);
   U667 : AOI221 port map( A => n247, B => U2_x_29_0_port, C => n262, D => 
                           U2_x_28_0_port, Q => U2_n333);
   U668 : INV3 port map( A => U2_n334, Q => U2_n249);
   U669 : AOI221 port map( A => n247, B => U2_x_30_7_port, C => n249, D => 
                           U2_x_29_7_port, Q => U2_n334);
   U670 : INV3 port map( A => U2_n335, Q => U2_n250);
   U671 : AOI221 port map( A => n248, B => U2_x_30_6_port, C => n261, D => 
                           U2_x_29_6_port, Q => U2_n335);
   U672 : INV3 port map( A => U2_n336, Q => U2_n251);
   U673 : AOI221 port map( A => n248, B => U2_x_30_5_port, C => n262, D => 
                           U2_x_29_5_port, Q => U2_n336);
   U674 : INV3 port map( A => U2_n337, Q => U2_n252);
   U675 : AOI221 port map( A => n248, B => U2_x_30_4_port, C => n261, D => 
                           U2_x_29_4_port, Q => U2_n337);
   U676 : INV3 port map( A => U2_n338, Q => U2_n253);
   U677 : AOI221 port map( A => n248, B => U2_x_30_3_port, C => n261, D => 
                           U2_x_29_3_port, Q => U2_n338);
   U678 : INV3 port map( A => U2_n339, Q => U2_n254);
   U679 : AOI221 port map( A => n248, B => U2_x_30_2_port, C => n249, D => 
                           U2_x_29_2_port, Q => U2_n339);
   U680 : INV3 port map( A => U2_n340, Q => U2_n255);
   U681 : AOI221 port map( A => n248, B => U2_x_30_1_port, C => n250, D => 
                           U2_x_29_1_port, Q => U2_n340);
   U682 : INV3 port map( A => U2_n341, Q => U2_n256);
   U683 : AOI221 port map( A => n248, B => U2_x_30_0_port, C => n261, D => 
                           U2_x_29_0_port, Q => U2_n341);
   U684 : INV3 port map( A => U2_n310, Q => U2_n257);
   U685 : AOI221 port map( A => n246, B => U2_x_31_7_port, C => n262, D => 
                           U2_x_30_7_port, Q => U2_n310);
   U686 : INV3 port map( A => U2_n311, Q => U2_n258);
   U687 : AOI221 port map( A => n246, B => U2_x_31_6_port, C => n262, D => 
                           U2_x_30_6_port, Q => U2_n311);
   U688 : INV3 port map( A => U2_n312, Q => U2_n259);
   U689 : AOI221 port map( A => n246, B => U2_x_31_5_port, C => n262, D => 
                           U2_x_30_5_port, Q => U2_n312);
   U690 : INV3 port map( A => U2_n313, Q => U2_n260);
   U691 : AOI221 port map( A => n246, B => U2_x_31_4_port, C => n250, D => 
                           U2_x_30_4_port, Q => U2_n313);
   U692 : INV3 port map( A => U2_n314, Q => U2_n261);
   U693 : AOI221 port map( A => n246, B => U2_x_31_3_port, C => n250, D => 
                           U2_x_30_3_port, Q => U2_n314);
   U694 : INV3 port map( A => U2_n315, Q => U2_n262);
   U695 : AOI221 port map( A => n247, B => U2_x_31_2_port, C => n262, D => 
                           U2_x_30_2_port, Q => U2_n315);
   U696 : INV3 port map( A => U2_n316, Q => U2_n263);
   U697 : AOI221 port map( A => n247, B => U2_x_31_1_port, C => n262, D => 
                           U2_x_30_1_port, Q => U2_n316);
   U698 : INV3 port map( A => U2_n317, Q => U2_n264);
   U699 : AOI221 port map( A => n247, B => U2_x_31_0_port, C => n250, D => 
                           U2_x_30_0_port, Q => U2_n317);
   U700 : NOR31 port map( A => n121, B => U6_n33, C => n19, Q => U6_n27);
   U701 : NAND22 port map( A => U7_n9, B => n148, Q => U7_n12);
   U702 : NAND22 port map( A => Filter_In(7), B => U9_n3, Q => U9_n10);
   U703 : NAND22 port map( A => Filter_In(6), B => U9_n3, Q => U9_n9);
   U704 : NAND22 port map( A => Filter_In(5), B => U9_n3, Q => U9_n8);
   U705 : NAND22 port map( A => Filter_In(4), B => U9_n3, Q => U9_n7);
   U706 : NAND22 port map( A => Filter_In(3), B => U9_n3, Q => U9_n6);
   U707 : NAND22 port map( A => Filter_In(2), B => U9_n3, Q => U9_n5);
   U708 : NAND22 port map( A => Filter_In(1), B => U9_n3, Q => U9_n4);
   U709 : NAND22 port map( A => Filter_In(0), B => U9_n3, Q => U9_n2);
   U710 : NAND22 port map( A => Accu_out_19_port, B => U5_n3, Q => U5_n10);
   U711 : NAND22 port map( A => Accu_out_18_port, B => U5_n3, Q => U5_n9);
   U712 : NAND22 port map( A => Accu_out_17_port, B => U5_n3, Q => U5_n8);
   U713 : NAND22 port map( A => Accu_out_16_port, B => U5_n3, Q => U5_n7);
   U714 : NAND22 port map( A => Accu_out_15_port, B => U5_n3, Q => U5_n6);
   U715 : NAND22 port map( A => Accu_out_14_port, B => U5_n3, Q => U5_n5);
   U716 : NAND22 port map( A => Accu_out_13_port, B => U5_n3, Q => U5_n4);
   U717 : NAND22 port map( A => Accu_out_12_port, B => U5_n3, Q => U5_n2);
   U718 : NAND22 port map( A => Accu_out_19_port, B => U6_n24, Q => 
                           U4_mult_add_27_aco_PROD_not_19_port);
   U719 : INV3 port map( A => U6_n25, Q => U6_n10);
   U720 : AOI2111 port map( A => U6_n26, B => U6_n11, C => Buff_OE, D => 
                           ack_F2ADC, Q => U6_n25);
   U721 : NAND31 port map( A => U6_n47, B => U6_n27, C => U6_n48, Q => U6_n26);
   U722 : AOI211 port map( A => n150, B => U7_n2, C => n56, Q => ADC_Rdb_port);
   U723 : NOR31 port map( A => n148, B => U7_n9, C => n56, Q => U7_n13);
   U724 : NOR31 port map( A => U8_n5, B => U8_pre_req_F2DAC, C => 
                           U8_current_state, Q => U8_N5_port);
   U725 : NOR21 port map( A => n56, B => U7_n10, Q => U7_n15);
   U726 : NOR21 port map( A => ADC_Eocb, B => n150, Q => U7_n11);
   U727 : INV3 port map( A => RESET, Q => n263);
   U728 : LOGIC0 port map( Q => LDACb);
   U729 : LOGIC1 port map( Q => CLRb);

end SYN_A;
