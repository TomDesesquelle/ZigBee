/softl1/AMS_410_ISR15/cds/HK_C35/LEF/c35b4/IOLIB_4M.lef