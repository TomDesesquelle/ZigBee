#  Last Change on: Fri Jul 06 13:37:13 2007
#  Owner: austriamicrosystems
#  Hit-Kit: Digital
#******
#  LEF Techfile created by ams_tech
#  
#  Process: C35B4
#  
#  TIPS-Document 
#         Nr.: ENG-182   Rev.: 3.0
#  DesignRules-Document 
#         Nr.: ENG-183   Rev.: 4.0
# 
#******

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 1000  ;
END UNITS

MANUFACTURINGGRID 0.025 ;

# Multiplication factor for CAP-Values is: 3.14

ANTENNAOUTPUTDIFFAREA 100000 ;
ANTENNAINOUTDIFFAREA 100000 ;

LAYER POLY1
  TYPE  MASTERSLICE ;
END POLY1

LAYER POLY2
  TYPE  MASTERSLICE ;
END POLY2

LAYER MET1
    TYPE ROUTING ;
    WIDTH 0.5 ;
    SPACING 0.45 ;
    SPACING 0.8 RANGE 10 10000 ;
    PITCH 1.3 ;
    OFFSET 0 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.000119 ;
    RESISTANCE RPERSQ 0.120000 ;
    EDGECAPACITANCE 0.000154 ;
    THICKNESS 0.665000 ;
    ANTENNASIDEAREARATIO 400 ;
END MET1

LAYER VIA1
    TYPE CUT ;
END VIA1
 
LAYER MET2
    TYPE ROUTING ;
    WIDTH 0.6 ;
    SPACING 0.5 ;
    SPACING 0.8 RANGE 10 10000 ;
    PITCH 1.4 ;
    OFFSET 0.7 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.000053 ;
    RESISTANCE RPERSQ 0.120000 ;
    EDGECAPACITANCE 0.000122 ;
    THICKNESS 0.640000 ;
    ANTENNASIDEAREARATIO 400 ;
END MET2
 
LAYER VIA2
    TYPE CUT ;
END VIA2
 
LAYER MET3
    TYPE ROUTING ;
    WIDTH 0.6 ;
    SPACING 0.5 ;
    SPACING 0.8 RANGE 10 10000 ;
    PITCH 1.3 ;
    OFFSET 0 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.000035 ;
    RESISTANCE RPERSQ 0.120000 ;
    EDGECAPACITANCE 0.000107 ;
    THICKNESS 0.640000 ;
    ANTENNASIDEAREARATIO 400 ;
END MET3
 
LAYER VIA3
    TYPE CUT ;
END VIA3
 
LAYER MET4
    TYPE ROUTING ;
    WIDTH 0.6 ;
    SPACING 0.6 ;
    SPACING 0.8 RANGE 10 10000 ;
    PITCH 1.4 ;
    OFFSET 0.7 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.000025 ;
    RESISTANCE RPERSQ 0.100000 ;
    EDGECAPACITANCE 0.000100 ;
    THICKNESS 0.925000 ;
    ANTENNASIDEAREARATIO 400 ;
END MET4


LAYER OVERLAP
    TYPE OVERLAP ;
END OVERLAP


# Via Met1-Met2 for normal routing
VIA VIA1_PR DEFAULT
    RESISTANCE 3 ;
    FOREIGN VIA1_C ;
    LAYER MET1 ;
        RECT -0.300000 -0.300000 0.300000 0.300000 ;
    LAYER VIA1 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
    LAYER MET2 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
END VIA1_PR

# Via Met2-Met3 for normal routing
VIA VIA2_PR DEFAULT
    RESISTANCE 3 ;
    FOREIGN VIA2_C ;
    LAYER MET2 ;
        RECT -0.300000 -0.300000 0.300000 0.300000 ;
    LAYER VIA2 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
    LAYER MET3 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
END VIA2_PR

# Via Met3-Met4 for normal routing
VIA VIA3_PR DEFAULT
    RESISTANCE 3 ;
    FOREIGN VIA3_C ;
    LAYER MET3 ;
        RECT -0.300000 -0.300000 0.300000 0.300000 ;
    LAYER VIA3 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
    LAYER MET4 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
END VIA3_PR

# Rule Via (needed for DEF import to DFII)
#VIA ruleVia
#        RESISTANCE 3 ;
#        LAYER MET1 ;
#          RECT -0.925000 -0.450000 0.925000 0.450000 ;
#        LAYER VIA1 ;
#          RECT -0.725000 -0.250000 -0.225000 0.250000 ;
#          RECT 0.225000 -0.250000 0.725000 0.250000 ;
#        LAYER MET2 ;
#          RECT -0.875000 -0.400000 0.875000 0.400000 ;
#END ruleVia
#
## Rule Via (needed for DEF import to DFII)
#VIA ruleVia2
#        RESISTANCE 3 ;
#        LAYER MET2 ;
#          RECT -0.925000 -0.450000 0.925000 0.450000 ;
#        LAYER VIA2 ;
#          RECT -0.725000 -0.250000 -0.225000 0.250000 ;
#          RECT 0.225000 -0.250000 0.725000 0.250000 ;
#        LAYER MET3 ;
#          RECT -0.875000 -0.400000 0.875000 0.400000 ;
#END ruleVia2
#
## Rule Via (needed for DEF import to DFII)
#VIA ruleVia3
#        RESISTANCE 3 ;
#        LAYER MET3 ;
#          RECT -0.925000 -0.450000 0.925000 0.450000 ;
#        LAYER VIA3 ;
#          RECT -0.725000 -0.250000 -0.225000 0.250000 ;
#          RECT 0.225000 -0.250000 0.725000 0.250000 ;
#        LAYER MET4 ;
#          RECT -0.875000 -0.400000 0.875000 0.400000 ;
#END ruleVia3
#
# Via Array for Wide-Met1/Wide-Met2
VIARULE VIA1W2W_G GENERATE
    LAYER MET2 ;
       DIRECTION VERTICAL ; 
       WIDTH 10 TO 1000.0 ; 
       OVERHANG 0.2 ;
       METALOVERHANG 0.00 ;

    LAYER MET1 ;
        DIRECTION HORIZONTAL ; 
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;

    LAYER VIA1 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.450000 BY 0.450000 ;
    RESISTANCE 3 ;
END VIA1W2W_G

# Via Array for Wide-Met1/Met2
# normal routing direction Met1 horizontal/Met2 vertical 
VIARULE VIA1W2_G GENERATE
    LAYER MET2 ;
        DIRECTION VERTICAL ; 
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;

    LAYER MET1 ;
        DIRECTION HORIZONTAL ; 
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;

    LAYER VIA1 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.450000 BY 0.450000 ;
    RESISTANCE 3 ;
END VIA1W2_G

# Via Array for Met1/Wide-Met2
# Normal routing direction Met1 horizontal / Met2 vertical
VIARULE VIA12W_G GENERATE
    LAYER MET2 ;
        DIRECTION VERTICAL ; 
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;

    LAYER MET1 ;
        DIRECTION HORIZONTAL ; 
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;

    LAYER VIA1 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.450 BY 0.450000 ;
    RESISTANCE 3 ;
END VIA12W_G

# Via Array for Wide-Met2/Wide-Met3
VIARULE VIA2W3W_G GENERATE
    LAYER MET2 ;
        DIRECTION HORIZONTAL ;
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;
 
    LAYER MET3 ;
        DIRECTION VERTICAL ;
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;
 
    LAYER VIA2 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.450000 BY 0.450000 ;
    RESISTANCE 3 ;
END VIA2W3W_G
 
# Via Array for Met2/Wide-Met3
# Normal routing direction Met2 vertical / Met3 horizontal
VIARULE VIA23W_G GENERATE
    LAYER MET2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;
 
    LAYER MET3 ;
        DIRECTION HORIZONTAL ;
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;
 
    LAYER VIA2 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.450000 BY 0.450000 ;
    RESISTANCE 3 ;
END VIA23W_G
 
# Via Array for Wide-Met2/Met3
# Normal routing direction Met2 vertical / Met3 horizontal
VIARULE VIA2W3_G GENERATE
    LAYER MET2 ;
        DIRECTION VERTICAL ;
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;
 
    LAYER MET3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.2 ; 
        METALOVERHANG 0.00 ;
 
    LAYER VIA2 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.450000 BY 0.450000 ;
    RESISTANCE 3 ;
END VIA2W3_G
 
# Via Array for Wide-Met3/Wide-Met4
VIARULE VIA3W4W_G GENERATE
    LAYER MET3 ;
        DIRECTION HORIZONTAL ;
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;
 
    LAYER MET4 ;
        DIRECTION VERTICAL ;
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;
 
    LAYER VIA3 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.450000 BY 0.450000 ;
    RESISTANCE 3 ;
END VIA3W4W_G
 
# Via Array for Met3/Wide-Met4
# Normal routing direction Met3 vertical / Met4 horizontal
VIARULE VIA34W_G GENERATE
    LAYER MET3 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;
 
    LAYER MET4 ;
        DIRECTION HORIZONTAL ;
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;
 
    LAYER VIA3 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.450000 BY 0.450000 ;
    RESISTANCE 3 ;
END VIA34W_G
 
# Via Array for Wide-Met3/Met4
# Normal routing direction Met3 vertical / Met4 horizontal
VIARULE VIA3W4_G GENERATE
    LAYER MET3 ;
        DIRECTION VERTICAL ;
        WIDTH 10 TO 1000.0 ; 
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;
 
    LAYER MET4 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.2 ; 
        METALOVERHANG 0.00 ;
 
    LAYER VIA3 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.450000 BY 0.450000 ;
    RESISTANCE 3 ;
END VIA3W4_G
 
# Via Array for Met1/Met2
VIARULE VIA12_G GENERATE
    LAYER MET2 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;

    LAYER MET1 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;

    LAYER VIA1 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.450000 BY 0.450000 ;
    RESISTANCE 3 ;
END VIA12_G

# Via Array for Met2/Met3
VIARULE VIA23_G GENERATE
    LAYER MET2 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;
 
    LAYER MET3 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;
 
    LAYER VIA2 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.450000 BY 0.450000 ;
    RESISTANCE 3 ;
END VIA23_G

# Via Array for Met3/Met4
VIARULE VIA34_G GENERATE
    LAYER MET3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;
 
    LAYER MET4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.2 ;
        METALOVERHANG 0.00 ;
 
    LAYER VIA3 ;
        RECT -0.250000 -0.250000 0.250000 0.250000 ;
        SPACING 0.450000 BY 0.450000 ;
    RESISTANCE 3 ;
END VIA34_G

SPACING
    SAMENET VIA1 VIA1 0.45 STACK ;
    SAMENET VIA2 VIA2 0.45 ;
    SAMENET VIA1 VIA2 0 STACK ;
    SAMENET VIA3 VIA3 0.45 ;
    SAMENET VIA2 VIA3 0 STACK ;
    SAMENET MET1 MET1 0.45 ;
    SAMENET MET2 MET2 0.5 STACK ;
    SAMENET MET3 MET3 0.5 STACK ;
    SAMENET MET4 MET4 0.6 STACK ;
END SPACING
 
SITE standard
    SYMMETRY y ;
    CLASS CORE ;
    SIZE 1.40 BY 13.00 ;
END standard

SITE portCellSite
    CLASS PAD ;
    SIZE 0.6 BY 0.6 ;
END portCellSite

SITE blockSite
    CLASS CORE  ;
    SIZE 1.00 BY 1.00 ;
END blockSite

SITE ioSite_P
    SYMMETRY y  ;
    CLASS pad  ;
    SIZE 0.10 BY 340.40 ;
END ioSite_P

SITE corner_P
    SYMMETRY x y r90 ;
    CLASS PAD ;
    SIZE 340.40 BY 340.40 ;
END corner_P


END LIBRARY
