`include ""

module msk_modulator_io2( 
